magic
tech sky130A
magscale 1 2
timestamp 1747754763
<< locali >>
rect 1487 621 3461 716
rect 395 367 479 563
rect 395 226 575 367
rect 395 -189 444 226
rect 483 -189 575 226
rect 395 -208 575 -189
rect 395 -564 479 -208
rect 395 -705 571 -564
rect 395 -1120 448 -705
rect 487 -1120 571 -705
rect 395 -1139 571 -1120
rect 395 -1334 479 -1139
rect 923 -1334 1007 563
rect 1483 -368 3457 -273
rect 1485 -693 3459 -598
rect 1489 -1683 3463 -1588
rect 395 -2454 479 -1704
rect 923 -1890 1007 -1704
rect 830 -2271 847 -1897
rect 923 -2258 940 -1890
rect 978 -2258 1007 -1890
rect 1048 -2024 3943 -1935
rect 923 -2454 1007 -2258
rect 1449 -2512 1558 -2024
rect 1044 -2602 1561 -2512
rect 3348 -2602 3506 -2024
rect 3796 -2598 3931 -2218
rect 1044 -2616 3506 -2602
rect 1044 -2676 3504 -2616
rect 1044 -2727 1063 -2676
rect 3409 -2727 3504 -2676
rect 1044 -2746 3504 -2727
rect 3326 -2816 3504 -2746
<< viali >>
rect 444 -189 483 226
rect 448 -1120 487 -705
rect 1446 264 1518 459
rect 3426 265 3498 460
rect 1455 -1041 1527 -846
rect 3426 -1041 3498 -846
rect 940 -2258 978 -1890
rect 1063 -2727 3409 -2676
<< metal1 >>
rect 978 568 1178 724
rect 677 524 1178 568
rect 1257 678 1457 727
rect 1257 629 2744 678
rect 1257 527 1457 629
rect 1724 542 1773 629
rect 677 519 1101 524
rect 438 226 490 236
rect 438 -189 444 226
rect 483 -189 490 226
rect 438 -199 490 -189
rect 441 -705 493 -696
rect 441 -1120 448 -705
rect 487 -1120 493 -705
rect 441 -1131 493 -1120
rect 677 -1228 726 519
rect 1719 518 1773 542
rect 1434 459 1531 469
rect 1434 264 1446 459
rect 1518 264 1531 459
rect 1434 251 1531 264
rect 1320 83 1387 99
rect 1320 -142 1387 -110
rect 1110 -209 1387 -142
rect 1110 -1796 1177 -209
rect 683 -1842 1177 -1796
rect 529 -2110 576 -1886
rect 300 -2310 576 -2110
rect 529 -2407 576 -2310
rect 683 -2348 717 -1842
rect 838 -1878 918 -1877
rect 838 -1890 991 -1878
rect 838 -2258 940 -1890
rect 978 -2258 991 -1890
rect 1110 -1979 1177 -1842
rect 1326 -1242 1393 -363
rect 1719 -647 1768 518
rect 2207 -261 2256 542
rect 2695 -200 2744 629
rect 3183 -131 3232 542
rect 3415 460 3509 472
rect 3415 265 3426 460
rect 3498 265 3509 460
rect 3415 253 3509 265
rect 3181 -200 3232 -131
rect 3181 -261 3230 -200
rect 2207 -310 3230 -261
rect 1719 -696 2744 -647
rect 1443 -846 1540 -836
rect 1443 -1041 1455 -846
rect 1527 -1041 1540 -846
rect 1443 -1054 1540 -1041
rect 1326 -1853 1393 -1435
rect 1719 -1790 1768 -696
rect 2207 -1576 2256 -768
rect 2695 -1510 2744 -696
rect 3183 -1484 3232 -768
rect 3414 -846 3511 -836
rect 3414 -1041 3426 -846
rect 3498 -1041 3511 -846
rect 3414 -1054 3511 -1041
rect 3181 -1510 3232 -1484
rect 3181 -1576 3230 -1510
rect 2117 -1624 3230 -1576
rect 2117 -1625 2641 -1624
rect 2714 -1625 3230 -1624
rect 1326 -1920 2597 -1853
rect 1110 -2046 1707 -1979
rect 1110 -2114 1177 -2046
rect 1110 -2148 1271 -2114
rect 838 -2269 991 -2258
rect 931 -2280 991 -2269
rect 1132 -2407 1179 -2194
rect 529 -2454 1179 -2407
rect 1237 -2431 1271 -2148
rect 1640 -2414 1707 -2046
rect 1763 -2154 1797 -2071
rect 2217 -2146 2247 -1920
rect 1767 -2158 1796 -2154
rect 1767 -2161 1802 -2158
rect 2215 -2159 2247 -2146
rect 1767 -2457 1796 -2161
rect 1866 -2368 2149 -2267
rect 2215 -2457 2244 -2159
rect 2530 -2406 2597 -1920
rect 2659 -2180 2695 -2055
rect 3105 -2146 3134 -1625
rect 3105 -2159 3140 -2146
rect 2667 -2185 2695 -2180
rect 2207 -2463 2244 -2457
rect 2663 -2464 2692 -2185
rect 2747 -2368 3030 -2267
rect 2660 -2474 2693 -2464
rect 3111 -2478 3140 -2159
rect 1044 -2672 3434 -2650
rect 3700 -2671 3734 -1781
rect 1044 -2727 1063 -2672
rect 3409 -2727 3434 -2672
rect 1044 -2746 3434 -2727
<< via1 >>
rect 1449 266 1517 458
rect 1320 -110 1387 83
rect 3428 265 3496 457
rect 1458 -1035 1526 -847
rect 1326 -1435 1393 -1242
rect 3429 -1039 3497 -847
rect 1063 -2676 3409 -2672
rect 1063 -2727 3409 -2676
<< metal2 >>
rect 428 -1161 657 739
rect 489 -1162 657 -1161
rect 778 266 1449 458
rect 1517 457 3490 458
rect 1517 266 3428 457
rect 778 265 3428 266
rect 3496 265 3504 457
rect 778 -430 937 265
rect 1300 -110 1320 83
rect 1387 -110 3488 83
rect 1331 -315 2282 -256
rect 1331 -391 1390 -315
rect 778 -839 928 -430
rect 778 -847 1244 -839
rect 778 -1035 1458 -847
rect 1526 -1035 3429 -847
rect 778 -1039 3429 -1035
rect 3497 -1039 3529 -847
rect 778 -1040 3529 -1039
rect 778 -1179 928 -1040
rect 780 -2500 928 -1179
rect 1312 -1435 1326 -1242
rect 1393 -1435 3485 -1242
rect 1149 -1628 2252 -1569
rect 1686 -1785 3548 -1742
rect 3857 -1846 4057 -1819
rect 2433 -1881 4057 -1846
rect 2433 -2036 2468 -1881
rect 3857 -1913 4057 -1881
rect 1919 -2071 2468 -2036
rect 2822 -2039 3578 -2038
rect 3857 -2039 4057 -2016
rect 2822 -2075 4057 -2039
rect 3541 -2076 4057 -2075
rect 3857 -2128 4057 -2076
rect 1305 -2600 1415 -2176
rect 1568 -2406 3671 -2203
rect 740 -2672 3970 -2600
rect 740 -2727 1063 -2672
rect 3409 -2727 3970 -2672
rect 740 -2800 3970 -2727
use pa_via  pa_via_0
timestamp 1717165164
transform 1 0 799 0 1 -4742
box -10 3586 63 4043
use pa_via  pa_via_1
timestamp 1717165164
transform 1 0 441 0 1 -4728
box -10 3586 63 4043
use pa_via  pa_via_2
timestamp 1717165164
transform 1 0 542 0 1 -4592
box -10 3586 63 4043
use pa_via  pa_via_3
timestamp 1717165164
transform 1 0 797 0 1 -3806
box -10 3586 63 4043
use pa_via  pa_via_4
timestamp 1717165164
transform 1 0 3805 0 1 -6252
box -10 3586 63 4043
use pa_via  pa_via_5
timestamp 1717165164
transform 1 0 540 0 1 -3659
box -10 3586 63 4043
use pa_via  pa_via_6
timestamp 1717165164
transform 1 0 438 0 1 -3796
box -10 3586 63 4043
use pa_via_short  pa_via_short_0
timestamp 1717168741
transform 1 0 -3624 0 1 -489
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_1
timestamp 1717168741
transform 1 0 -4131 0 1 -291
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_2
timestamp 1717168741
transform 1 0 -3106 0 1 1773
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_3
timestamp 1717168741
transform 1 0 -3381 0 1 2140
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_4
timestamp 1717168741
transform 1 0 -2890 0 1 2154
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_5
timestamp 1717168741
transform 1 0 -2399 0 1 2148
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_6
timestamp 1717168741
transform 1 0 -1914 0 1 2148
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_7
timestamp 1717168741
transform 1 0 -2612 0 1 1781
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_8
timestamp 1717168741
transform 1 0 -2142 0 1 1767
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_9
timestamp 1717168741
transform 1 0 -2887 0 1 844
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_10
timestamp 1717168741
transform 1 0 -1657 0 1 1770
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_11
timestamp 1717168741
transform 1 0 -1657 0 1 448
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_12
timestamp 1717168741
transform 1 0 -2139 0 1 454
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_13
timestamp 1717168741
transform 1 0 -2627 0 1 451
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_14
timestamp 1717168741
transform 1 0 -3106 0 1 454
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_15
timestamp 1717168741
transform 1 0 -3360 0 1 846
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_16
timestamp 1717168741
transform 1 0 -2396 0 1 855
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_17
timestamp 1717168741
transform 1 0 -1916 0 1 844
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_18
timestamp 1717168741
transform 1 0 -2648 0 1 -522
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_19
timestamp 1717168741
transform 1 0 -1348 0 1 -520
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_20
timestamp 1717168741
transform 1 0 -1759 0 1 -520
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_22
timestamp 1717168741
transform 1 0 -3834 0 1 195
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_24
timestamp 1717168741
transform 1 0 -3618 0 1 1322
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_25
timestamp 1717168741
transform 0 1 4006 -1 0 3380
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_26
timestamp 1717168741
transform 0 1 4091 -1 0 4693
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_28
timestamp 1717168741
transform 0 1 3541 -1 0 3218
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_29
timestamp 1717168741
transform 0 1 3639 -1 0 2918
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_30
timestamp 1717168741
transform 0 1 4529 -1 0 2919
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_32
timestamp 1717168741
transform 0 1 5426 -1 0 3220
box 4944 -1889 5010 -1683
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_0 paramcells
timestamp 1717168741
transform 1 0 1741 0 1 -1140
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_1
timestamp 1717168741
transform 1 0 2227 0 1 -1140
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_2
timestamp 1717168741
transform 1 0 2713 0 1 -1140
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_3
timestamp 1717168741
transform 1 0 3199 0 1 -1140
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_4
timestamp 1717168741
transform 1 0 701 0 1 80
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  sky130_fd_pr__pfet_01v8_hvt_3HBZVM_5
timestamp 1717168741
transform 1 0 701 0 1 -852
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  XM1
timestamp 1717168741
transform 1 0 3201 0 1 170
box -296 -519 296 519
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM2 paramcells
timestamp 1717168741
transform 1 0 1782 0 1 -2317
box -288 -358 288 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM3
timestamp 1717168741
transform 1 0 2228 0 1 -2317
box -288 -358 288 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM4
timestamp 1717168741
transform 1 0 2674 0 1 -2317
box -288 -358 288 358
use sky130_fd_pr__nfet_03v3_nvt_UNEQ2N  XM5
timestamp 1717168741
transform 1 0 3120 0 1 -2317
box -288 -358 288 358
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  XM10
timestamp 1717168741
transform 1 0 1743 0 1 170
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  XM11
timestamp 1717168741
transform 1 0 2229 0 1 170
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_hvt_3HBZVM  XM12
timestamp 1717168741
transform 1 0 2715 0 1 170
box -296 -519 296 519
use sky130_fd_pr__nfet_03v3_nvt_WSEQJ8  XM15 paramcells
timestamp 1717166647
transform 1 0 3720 0 1 -2409
box -278 -458 278 458
use sky130_fd_pr__nfet_01v8_PVEW3M  XM18 paramcells
timestamp 1717166647
transform 1 0 1258 0 1 -2279
box -246 -310 246 310
use sky130_fd_pr__pfet_01v8_3HY9VM  XM19 paramcells
timestamp 1717166647
transform 1 0 701 0 1 -2084
box -296 -419 296 419
<< labels >>
flabel metal2 740 -2800 940 -2600 0 FreeSans 256 0 0 0 dvss
port 7 nsew
flabel metal2 1044 -1039 1244 -839 0 FreeSans 256 0 0 0 dvddb
port 2 nsew
flabel metal1 1257 527 1457 727 0 FreeSans 256 0 0 0 clkb
port 3 nsew
flabel metal2 431 539 631 739 0 FreeSans 256 0 0 0 dvdd
port 0 nsew
flabel metal1 300 -2310 500 -2110 0 FreeSans 256 0 0 0 vout
port 4 nsew
flabel metal1 978 524 1178 724 0 FreeSans 256 0 0 0 enab
port 1 nsew
flabel metal2 3857 -1913 4057 -1819 0 FreeSans 256 0 0 0 opos
port 6 nsew
flabel metal2 3857 -2128 4057 -2016 0 FreeSans 256 0 0 0 oneg
port 5 nsew
<< end >>
