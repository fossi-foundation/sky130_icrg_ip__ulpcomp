magic
tech sky130A
magscale 1 2
timestamp 1718247345
<< dnwell >>
rect 402 -4779 4688 -2850
<< nwell >>
rect 293 -3056 4797 -2727
rect 293 -4573 608 -3056
rect 2297 -4573 2865 -3056
rect 4482 -4573 4797 -3056
rect 293 -4888 4797 -4573
<< mvpsubdiff >>
rect 5434 2864 5494 2898
rect 7903 2864 7963 2898
rect 5434 2838 5468 2864
rect 5434 -538 5468 -512
rect 7929 2838 7963 2864
rect 7929 -538 7963 -512
rect 5434 -572 5494 -538
rect 7903 -572 7963 -538
<< mvnsubdiff >>
rect 359 -2833 4731 -2807
rect 359 -2854 456 -2833
rect 359 -4742 379 -2854
rect 413 -2869 456 -2854
rect 4616 -2869 4731 -2833
rect 413 -2881 4731 -2869
rect 413 -4742 433 -2881
rect 359 -4748 433 -4742
rect 4657 -2919 4731 -2881
rect 4657 -4742 4677 -2919
rect 4711 -4742 4731 -2919
rect 4657 -4748 4731 -4742
rect 359 -4768 4731 -4748
rect 359 -4802 439 -4768
rect 4651 -4802 4731 -4768
rect 359 -4822 4731 -4802
<< mvpsubdiffcont >>
rect 5494 2864 7903 2898
rect 5434 -512 5468 2838
rect 7929 -512 7963 2838
rect 5494 -572 7903 -538
<< mvnsubdiffcont >>
rect 379 -4742 413 -2854
rect 456 -2869 4616 -2833
rect 4677 -4742 4711 -2919
rect 439 -4802 4651 -4768
<< locali >>
rect 1887 4377 4796 4389
rect 1887 4340 1915 4377
rect 4724 4340 4796 4377
rect 1887 4317 4796 4340
rect 19 3148 160 4136
rect 1187 3146 1328 4134
rect 5434 2864 5494 2898
rect 7903 2864 7963 2898
rect 5434 2838 7963 2864
rect 22 1745 163 2733
rect 1190 1744 1331 2732
rect -6 1519 1347 1596
rect 1887 1560 4794 1583
rect 1887 1523 1923 1560
rect 4742 1523 4794 1560
rect 1887 1510 4794 1523
rect -3 908 1350 985
rect 1889 972 4788 982
rect 1889 926 1916 972
rect 4767 926 4788 972
rect 1889 917 4788 926
rect 21 -243 162 745
rect 1190 -238 1331 750
rect 5433 -512 5434 -459
rect 5468 2785 7929 2838
rect 5468 -459 5540 2785
rect 5640 2365 5745 2378
rect 5640 2158 5651 2365
rect 5732 2158 5745 2365
rect 5640 2145 5745 2158
rect 7270 1592 7472 1605
rect 7270 1486 7286 1592
rect 7458 1486 7472 1592
rect 7270 1471 7472 1486
rect 5641 734 5746 747
rect 5641 527 5652 734
rect 5733 527 5746 734
rect 5641 514 5746 527
rect 7270 -36 7472 -23
rect 7270 -142 7286 -36
rect 7458 -142 7472 -36
rect 7270 -157 7472 -142
rect 7858 -459 7929 2785
rect 5468 -512 7929 -459
rect 5433 -538 7963 -512
rect 5433 -567 5494 -538
rect 5434 -572 5494 -567
rect 7903 -572 7963 -538
rect 22 -1647 163 -659
rect 1188 -1647 1329 -659
rect -3 -1881 1350 -1804
rect 1882 -1819 4792 -1813
rect 1882 -1865 1916 -1819
rect 4767 -1865 4792 -1819
rect 1882 -1884 4792 -1865
rect 615 -2826 4711 -2811
rect 615 -2833 642 -2826
rect 379 -2854 456 -2833
rect 413 -2869 456 -2854
rect 4666 -2864 4711 -2826
rect 4616 -2869 4711 -2864
rect 615 -2880 4711 -2869
rect 4677 -2919 4711 -2880
rect 1119 -3091 2290 -3079
rect 1119 -3143 1153 -3091
rect 1119 -3163 2290 -3143
rect 1119 -3843 1178 -3163
rect 1119 -3852 1197 -3843
rect 1119 -4051 1133 -3852
rect 1185 -4051 1197 -3852
rect 1119 -4062 1197 -4051
rect 1119 -4457 1178 -4062
rect 1602 -4457 1772 -3163
rect 2201 -3846 2290 -3163
rect 2180 -3858 2290 -3846
rect 2180 -4051 2195 -3858
rect 2276 -4051 2290 -3858
rect 2180 -4061 2290 -4051
rect 2201 -4457 2290 -4061
rect 1119 -4473 2290 -4457
rect 1119 -4525 1163 -4473
rect 1119 -4541 2290 -4525
rect 2855 -3091 4041 -3079
rect 4009 -3143 4041 -3091
rect 2855 -3163 4041 -3143
rect 2855 -4112 2971 -3163
rect 2855 -4305 2867 -4112
rect 2968 -4305 2971 -4112
rect 2855 -4457 2971 -4305
rect 3394 -4457 3564 -3163
rect 3982 -4457 4041 -3163
rect 2855 -4473 4041 -4457
rect 4019 -4525 4041 -4473
rect 2855 -4541 4041 -4525
rect 379 -4746 413 -4742
rect 4677 -4746 4711 -4742
rect 371 -4763 4720 -4746
rect 371 -4804 388 -4763
rect 4681 -4804 4720 -4763
rect 371 -4821 4720 -4804
<< viali >>
rect 1915 4340 4724 4377
rect 1923 1523 4742 1560
rect 1916 926 4767 972
rect 5651 2158 5732 2365
rect 7286 1486 7458 1592
rect 5652 527 5733 734
rect 7286 -142 7458 -36
rect 1916 -1865 4767 -1819
rect 642 -2833 4666 -2826
rect 642 -2864 4616 -2833
rect 4616 -2864 4666 -2833
rect 1153 -3143 2290 -3091
rect 1133 -4051 1185 -3852
rect 2195 -4051 2276 -3858
rect 1163 -4525 2290 -4473
rect 2855 -3143 4009 -3091
rect 2867 -4305 2968 -4112
rect 2855 -4525 4019 -4473
rect 388 -4768 4681 -4763
rect 388 -4802 439 -4768
rect 439 -4802 4651 -4768
rect 4651 -4802 4681 -4768
rect 388 -4804 4681 -4802
<< metal1 >>
rect 1887 4377 5314 4388
rect 1887 4340 1915 4377
rect 4724 4340 5314 4377
rect 1887 4324 5314 4340
rect 1887 4317 4908 4324
rect 4885 4229 4908 4317
rect 5291 4229 5314 4324
rect -280 2971 -80 3055
rect 275 2971 322 4226
rect 533 2971 580 4226
rect 791 2971 838 4226
rect 1049 2971 1096 4226
rect -280 2923 1546 2971
rect 2157 2961 2204 4223
rect 2415 2961 2462 4223
rect 2673 2961 2720 4223
rect 2931 2961 2978 4223
rect 3189 2961 3236 4223
rect 3447 2961 3494 4223
rect 3705 2961 3752 4223
rect 3963 2961 4010 4223
rect 4221 2961 4268 4223
rect 4479 2961 4526 4223
rect 4885 4211 5314 4229
rect -280 2922 248 2923
rect -280 2855 -80 2922
rect 275 1733 322 2832
rect 533 1751 580 2832
rect 791 1786 838 2832
rect 271 1681 322 1733
rect 529 1681 580 1751
rect 787 1681 838 1786
rect 1049 1746 1096 2832
rect 1045 1681 1096 1746
rect -274 1380 -74 1437
rect 271 1380 318 1681
rect 529 1380 576 1681
rect 787 1380 834 1681
rect 1045 1380 1092 1681
rect -274 1332 1397 1380
rect -274 1237 -74 1332
rect 1484 1275 1546 2923
rect 2152 2919 4986 2961
rect 2157 1678 2204 2919
rect 2415 1678 2462 2919
rect 2673 1678 2720 2919
rect 2931 1678 2978 2919
rect 3189 1678 3236 2919
rect 3447 1678 3494 2919
rect 3705 1678 3752 2919
rect 3963 1678 4010 2919
rect 4221 1678 4268 2919
rect 4479 1678 4526 2919
rect 4944 2251 4986 2919
rect 5450 2795 7948 2899
rect 5450 2687 7130 2795
rect 7520 2687 7948 2795
rect 5450 2668 7948 2687
rect 5640 2365 5745 2378
rect 5640 2251 5651 2365
rect 4944 2203 5651 2251
rect 5640 2158 5651 2203
rect 5732 2158 5745 2365
rect 5640 2145 5745 2158
rect 5661 1890 5867 2060
rect 6261 1890 7765 2060
rect 4885 1609 5314 1619
rect 4885 1581 4898 1609
rect 1887 1560 4898 1581
rect 1887 1523 1923 1560
rect 4742 1523 4898 1560
rect 1887 1510 4898 1523
rect 4885 1484 4898 1510
rect 5303 1484 5314 1609
rect 4885 1473 5314 1484
rect 7270 1592 7472 1605
rect 7270 1486 7286 1592
rect 7458 1569 7472 1592
rect 7642 1569 7842 1660
rect 7458 1513 7842 1569
rect 7458 1486 7472 1513
rect 7270 1471 7472 1486
rect 7642 1460 7842 1513
rect 271 1227 1546 1275
rect 271 -328 318 1227
rect 529 -328 576 1227
rect 787 -328 834 1227
rect 1045 -328 1092 1227
rect 5653 1076 7137 1246
rect 7511 1076 7757 1246
rect 1886 972 4834 1003
rect 1484 -435 1546 957
rect 1886 926 1916 972
rect 4767 926 4834 972
rect 1886 902 4834 926
rect 2153 -432 2200 813
rect 2411 -432 2458 813
rect 2669 -432 2716 813
rect 2927 -432 2974 813
rect 3185 -432 3232 813
rect 3443 -432 3490 813
rect 3701 -432 3748 813
rect 3959 -432 4006 813
rect 4217 -432 4264 813
rect 4475 -432 4522 813
rect 4742 220 4834 902
rect 5641 734 5746 747
rect 5641 653 5652 734
rect 4742 -217 4754 220
rect 4826 -217 4834 220
rect 4742 -227 4834 -217
rect 5294 605 5652 653
rect 5294 -216 5336 605
rect 5641 527 5652 605
rect 5733 527 5746 734
rect 5641 514 5746 527
rect 5659 258 5866 428
rect 6260 258 7763 428
rect 7270 -36 7472 -23
rect 7270 -142 7286 -36
rect 7458 -55 7472 -36
rect 7630 -55 7830 38
rect 7458 -111 7830 -55
rect 7458 -142 7472 -111
rect 7270 -157 7472 -142
rect 7630 -162 7830 -111
rect 5294 -432 5334 -216
rect 249 -468 1546 -435
rect 271 -1729 318 -468
rect 529 -1729 576 -468
rect 787 -1729 834 -468
rect 1045 -1729 1092 -468
rect 2146 -474 5352 -432
rect 5653 -471 7121 -370
rect 7519 -471 7765 -370
rect 5653 -474 7765 -471
rect 2153 -1732 2200 -474
rect 2411 -1732 2458 -474
rect 2669 -1732 2716 -474
rect 2927 -1732 2974 -474
rect 3185 -1732 3232 -474
rect 3443 -1732 3490 -474
rect 3701 -1732 3748 -474
rect 3959 -1732 4006 -474
rect 4217 -1732 4264 -474
rect 4475 -1732 4522 -474
rect 4739 -1186 4838 -1171
rect 4739 -1629 4747 -1186
rect 4829 -1629 4838 -1186
rect 4739 -1804 4838 -1629
rect 1870 -1819 4838 -1804
rect 1870 -1865 1916 -1819
rect 4767 -1865 4838 -1819
rect 1870 -1905 4838 -1865
rect 5294 -2024 5334 -474
rect 2640 -2064 5334 -2024
rect 4885 -2789 5314 -2778
rect 4885 -2813 4901 -2789
rect 615 -2826 4901 -2813
rect 615 -2864 642 -2826
rect 4666 -2864 4901 -2826
rect 615 -2880 4901 -2864
rect 4885 -2908 4901 -2880
rect 5299 -2908 5314 -2789
rect 4885 -2920 5314 -2908
rect 1121 -3091 2315 -3076
rect 1121 -3143 1153 -3091
rect 2290 -3143 2315 -3091
rect 1121 -3165 2315 -3143
rect 2550 -3212 2596 -2947
rect 2828 -3091 4040 -3076
rect 2828 -3143 2855 -3091
rect 4009 -3143 4040 -3091
rect 2828 -3156 2871 -3143
rect 3953 -3156 4040 -3143
rect 2828 -3165 4040 -3156
rect 1344 -3253 2596 -3212
rect 3128 -3253 3872 -3212
rect 1120 -3852 1197 -3843
rect 1120 -4051 1133 -3852
rect 1185 -4051 1197 -3852
rect 1120 -4062 1197 -4051
rect 1371 -4377 1408 -3256
rect 1965 -4379 2002 -3258
rect 3195 -3260 3280 -3253
rect 3787 -3258 3872 -3253
rect 3158 -3282 3280 -3260
rect 2180 -3858 2289 -3846
rect 2180 -4051 2195 -3858
rect 2276 -4051 2289 -3858
rect 2180 -4061 2289 -4051
rect 2855 -4112 2982 -4102
rect 2855 -4305 2867 -4112
rect 2968 -4305 2982 -4112
rect 2855 -4318 2982 -4305
rect 3158 -4381 3195 -3282
rect 3234 -3331 3280 -3282
rect 3752 -3282 3872 -3258
rect 3752 -4379 3789 -3282
rect 3826 -3321 3872 -3282
rect 1121 -4473 2315 -4457
rect 1121 -4525 1163 -4473
rect 2290 -4525 2315 -4473
rect 1121 -4541 2315 -4525
rect 2828 -4473 4043 -4457
rect 2828 -4525 2855 -4473
rect 4019 -4525 4043 -4473
rect 2828 -4541 4043 -4525
rect 4885 -4669 5314 -4653
rect 4885 -4746 4902 -4669
rect 371 -4763 4902 -4746
rect 371 -4804 388 -4763
rect 4681 -4804 4902 -4763
rect 371 -4805 4902 -4804
rect 5295 -4805 5314 -4669
rect 371 -4821 5314 -4805
<< via1 >>
rect 4908 4229 5291 4324
rect 7130 2687 7520 2795
rect 5867 1871 6261 2087
rect 6494 1769 6882 1826
rect 4898 1484 5303 1609
rect 7137 1072 7511 1257
rect 4754 -217 4826 220
rect 5866 244 6260 460
rect 6494 141 6882 198
rect 7121 -471 7519 -360
rect 4747 -1629 4829 -1186
rect 4901 -2908 5299 -2789
rect 2871 -3143 3953 -3091
rect 2871 -3156 3953 -3143
rect 1133 -4051 1185 -3852
rect 2195 -4051 2276 -3858
rect 2867 -4305 2968 -4112
rect 4902 -4805 5295 -4669
<< metal2 >>
rect 4885 4324 5314 4342
rect 4885 4229 4908 4324
rect 5291 4229 5314 4324
rect 4885 4211 5314 4229
rect 116 4106 1818 4115
rect 116 3674 982 4106
rect 1140 3674 1818 4106
rect 116 3656 1818 3674
rect 2018 4100 5315 4115
rect 2018 3668 2098 4100
rect 2252 3668 2614 4100
rect 2768 3668 3130 4100
rect 3284 3668 3646 4100
rect 3800 3668 4162 4100
rect 4316 4099 5315 4100
rect 4316 3668 4898 4099
rect 2018 3667 4898 3668
rect 5297 3667 5315 4099
rect 2018 3656 5315 3667
rect 116 3596 1816 3610
rect 116 3164 478 3596
rect 636 3164 1816 3596
rect 116 3151 1816 3164
rect 2011 3590 4680 3610
rect 2011 3169 2358 3590
rect 2511 3169 2874 3590
rect 3027 3169 3390 3590
rect 3543 3169 3906 3590
rect 4059 3169 4422 3590
rect 4575 3169 4680 3590
rect 2011 3151 4680 3169
rect 116 2719 1816 2722
rect 116 2287 729 2719
rect 887 2718 1816 2719
rect 2018 2721 5375 2722
rect 5849 2721 6284 2869
rect 887 2287 1818 2718
rect 116 2263 1818 2287
rect 2015 2261 2017 2718
rect 2018 2706 6284 2721
rect 2018 2704 4900 2706
rect 2018 2272 2098 2704
rect 2252 2272 2614 2704
rect 2768 2272 3130 2704
rect 3284 2272 3646 2704
rect 3800 2272 4162 2704
rect 4316 2279 4900 2704
rect 5295 2279 6284 2706
rect 4316 2272 6284 2279
rect 2018 2263 6284 2272
rect 4668 2262 6284 2263
rect 116 2209 1816 2215
rect 116 1777 224 2209
rect 382 1777 1816 2209
rect 2015 2194 4680 2215
rect 2015 2179 2358 2194
rect 116 1756 1816 1777
rect 2011 1773 2358 2179
rect 2511 1773 2874 2194
rect 3027 1773 3390 2194
rect 3543 1773 3906 2194
rect 4059 1773 4422 2194
rect 4575 1773 4680 2194
rect 2011 1756 4680 1773
rect 5849 2087 6284 2262
rect 5849 1871 5867 2087
rect 6261 1871 6284 2087
rect 4885 1609 5314 1619
rect 4885 1484 4898 1609
rect 5303 1484 5314 1609
rect 4885 1473 5314 1484
rect 1418 1325 1549 1391
rect 1482 998 1549 1325
rect 1485 997 1547 998
rect 116 720 4687 733
rect 116 288 979 720
rect 1137 717 4687 720
rect 1137 296 2101 717
rect 2254 296 3135 717
rect 3288 714 4687 717
rect 3288 296 4165 714
rect 1137 293 4165 296
rect 4318 293 4687 714
rect 1137 288 4687 293
rect 116 274 4687 288
rect 5849 460 6284 1871
rect 5849 244 5866 460
rect 6260 244 6284 460
rect 116 221 1818 229
rect 116 -211 474 221
rect 632 -211 1818 221
rect 116 -230 1818 -211
rect 2018 220 4835 229
rect 2018 208 4754 220
rect 2018 -213 2358 208
rect 2511 -213 2874 208
rect 3027 -213 3390 208
rect 3543 -213 3906 208
rect 4059 -213 4422 208
rect 4575 -213 4754 208
rect 2018 -217 4754 -213
rect 4826 -217 4835 220
rect 2018 -230 4835 -217
rect 5849 -581 6284 244
rect 6471 1826 6906 2870
rect 6471 1769 6494 1826
rect 6882 1769 6906 1826
rect 6471 198 6906 1769
rect 6471 141 6494 198
rect 6882 141 6906 198
rect 6471 -596 6906 141
rect 7105 2795 7540 2853
rect 7105 2687 7130 2795
rect 7520 2687 7540 2795
rect 7105 1257 7540 2687
rect 7105 1072 7137 1257
rect 7511 1072 7540 1257
rect 7105 -360 7540 1072
rect 7105 -471 7121 -360
rect 7519 -471 7540 -360
rect 7105 -566 7540 -471
rect 116 -686 4680 -673
rect 116 -688 3649 -686
rect 116 -1120 728 -688
rect 886 -698 3649 -688
rect 886 -1119 2615 -698
rect 2768 -1107 3649 -698
rect 3802 -1107 4680 -686
rect 2768 -1119 4680 -1107
rect 886 -1120 4680 -1119
rect 116 -1132 4680 -1120
rect 116 -1190 1818 -1177
rect 116 -1622 227 -1190
rect 385 -1622 1818 -1190
rect 116 -1636 1818 -1622
rect 2018 -1186 4840 -1177
rect 2018 -1188 4747 -1186
rect 2018 -1609 2358 -1188
rect 2511 -1609 2874 -1188
rect 3027 -1609 3390 -1188
rect 3543 -1609 3906 -1188
rect 4059 -1609 4422 -1188
rect 4575 -1609 4747 -1188
rect 2018 -1629 4747 -1609
rect 4829 -1629 4840 -1186
rect 2018 -1636 4840 -1629
rect 2541 -2968 2598 -2062
rect 4885 -2789 5314 -2778
rect 4885 -2908 4901 -2789
rect 5299 -2908 5314 -2789
rect 4885 -2920 5314 -2908
rect -303 -3087 4049 -3075
rect -303 -3233 -283 -3087
rect 105 -3091 4049 -3087
rect 105 -3156 2871 -3091
rect 3953 -3156 4049 -3091
rect 105 -3233 4049 -3156
rect -303 -3253 4049 -3233
rect 210 -3317 3892 -3308
rect 210 -3514 471 -3317
rect 636 -3338 3892 -3317
rect 5116 -3338 5316 -3233
rect 636 -3433 5316 -3338
rect 636 -3434 5116 -3433
rect 636 -3514 3892 -3434
rect 210 -3523 3892 -3514
rect 210 -3581 3897 -3570
rect 210 -3778 221 -3581
rect 386 -3589 3897 -3581
rect 5116 -3589 5316 -3505
rect 386 -3685 5316 -3589
rect 386 -3778 3897 -3685
rect 5116 -3705 5316 -3685
rect 210 -3785 3897 -3778
rect 1102 -3852 3893 -3846
rect 1102 -4051 1133 -3852
rect 1185 -3858 3893 -3852
rect 1185 -4051 2195 -3858
rect 2276 -4051 3893 -3858
rect 1102 -4062 3893 -4051
rect -305 -4111 3888 -4102
rect -305 -4309 -297 -4111
rect 112 -4112 3888 -4111
rect 112 -4305 2867 -4112
rect 2968 -4305 3888 -4112
rect 112 -4309 3888 -4305
rect -305 -4318 3888 -4309
rect 4885 -4669 5314 -4653
rect 4885 -4805 4902 -4669
rect 5295 -4805 5314 -4669
rect 4885 -4821 5314 -4805
<< via2 >>
rect 4908 4229 5291 4324
rect 982 3674 1140 4106
rect 2098 3668 2252 4100
rect 2614 3668 2768 4100
rect 3130 3668 3284 4100
rect 3646 3668 3800 4100
rect 4162 3668 4316 4100
rect 4898 3667 5297 4099
rect 478 3164 636 3596
rect 2358 3169 2511 3590
rect 2874 3169 3027 3590
rect 3390 3169 3543 3590
rect 3906 3169 4059 3590
rect 4422 3169 4575 3590
rect 729 2287 887 2719
rect 2098 2272 2252 2704
rect 2614 2272 2768 2704
rect 3130 2272 3284 2704
rect 3646 2272 3800 2704
rect 4162 2272 4316 2704
rect 4900 2279 5295 2706
rect 224 1777 382 2209
rect 2358 1773 2511 2194
rect 2874 1773 3027 2194
rect 3390 1773 3543 2194
rect 3906 1773 4059 2194
rect 4422 1773 4575 2194
rect 4898 1484 5303 1609
rect 979 288 1137 720
rect 2101 296 2254 717
rect 3135 296 3288 717
rect 4165 293 4318 714
rect 474 -211 632 221
rect 2358 -213 2511 208
rect 2874 -213 3027 208
rect 3390 -213 3543 208
rect 3906 -213 4059 208
rect 4422 -213 4575 208
rect 728 -1120 886 -688
rect 2615 -1119 2768 -698
rect 3649 -1107 3802 -686
rect 227 -1622 385 -1190
rect 2358 -1609 2511 -1188
rect 2874 -1609 3027 -1188
rect 3390 -1609 3543 -1188
rect 3906 -1609 4059 -1188
rect 4422 -1609 4575 -1188
rect 4901 -2908 5299 -2789
rect -283 -3233 105 -3087
rect 471 -3514 636 -3317
rect 221 -3778 386 -3581
rect -297 -4309 112 -4111
rect 4902 -4805 5295 -4669
<< metal3 >>
rect -305 -3075 124 4434
rect 4885 4324 5314 4550
rect 211 2209 398 4262
rect 211 1777 224 2209
rect 382 1777 398 2209
rect 211 -1190 398 1777
rect 211 -1622 227 -1190
rect 385 -1622 398 -1190
rect -305 -3087 125 -3075
rect -305 -3233 -283 -3087
rect 105 -3233 125 -3087
rect -305 -3253 125 -3233
rect -305 -4111 124 -3253
rect 211 -3581 398 -1622
rect 211 -3778 221 -3581
rect 386 -3778 398 -3581
rect 211 -3786 398 -3778
rect 463 3596 650 4262
rect 463 3164 478 3596
rect 636 3164 650 3596
rect 463 221 650 3164
rect 463 -211 474 221
rect 632 -211 650 221
rect 463 -3317 650 -211
rect 715 2719 902 4262
rect 715 2287 729 2719
rect 887 2287 902 2719
rect 715 -688 902 2287
rect 715 -1120 728 -688
rect 886 -1120 902 -688
rect 715 -1761 902 -1120
rect 967 4106 1154 4262
rect 967 3674 982 4106
rect 1140 3674 1154 4106
rect 967 720 1154 3674
rect 2083 4100 2271 4264
rect 2083 3668 2098 4100
rect 2252 3668 2271 4100
rect 2083 2704 2271 3668
rect 2083 2272 2098 2704
rect 2252 2272 2271 2704
rect 2083 1409 2271 2272
rect 2341 3590 2529 4264
rect 2341 3169 2358 3590
rect 2511 3169 2529 3590
rect 2341 2194 2529 3169
rect 2341 1773 2358 2194
rect 2511 1773 2529 2194
rect 967 288 979 720
rect 1137 288 1154 720
rect 967 -1761 1154 288
rect 2083 717 2271 1241
rect 2083 296 2101 717
rect 2254 296 2271 717
rect 2083 -1741 2271 296
rect 2341 208 2529 1773
rect 2599 4100 2787 4264
rect 2599 3668 2614 4100
rect 2768 3668 2787 4100
rect 2599 2704 2787 3668
rect 2599 2272 2614 2704
rect 2768 2272 2787 2704
rect 2599 1409 2787 2272
rect 2857 3590 3045 4264
rect 2857 3169 2874 3590
rect 3027 3169 3045 3590
rect 2857 2194 3045 3169
rect 2857 1773 2874 2194
rect 3027 1773 3045 2194
rect 2341 -213 2358 208
rect 2511 -213 2529 208
rect 2341 -1188 2529 -213
rect 2341 -1609 2358 -1188
rect 2511 -1609 2529 -1188
rect 2341 -1741 2529 -1609
rect 2599 -698 2787 1241
rect 2599 -1119 2615 -698
rect 2768 -1119 2787 -698
rect 2599 -1741 2787 -1119
rect 2857 208 3045 1773
rect 3115 4100 3303 4264
rect 3115 3668 3130 4100
rect 3284 3668 3303 4100
rect 3115 2704 3303 3668
rect 3115 2272 3130 2704
rect 3284 2272 3303 2704
rect 3115 1409 3303 2272
rect 3373 3590 3561 4264
rect 3373 3169 3390 3590
rect 3543 3169 3561 3590
rect 3373 2194 3561 3169
rect 3373 1773 3390 2194
rect 3543 1773 3561 2194
rect 2857 -213 2874 208
rect 3027 -213 3045 208
rect 2857 -1188 3045 -213
rect 2857 -1609 2874 -1188
rect 3027 -1609 3045 -1188
rect 2857 -1741 3045 -1609
rect 3115 717 3303 1241
rect 3115 296 3135 717
rect 3288 296 3303 717
rect 3115 -1741 3303 296
rect 3373 208 3561 1773
rect 3631 4100 3819 4264
rect 3631 3668 3646 4100
rect 3800 3668 3819 4100
rect 3631 2704 3819 3668
rect 3631 2272 3646 2704
rect 3800 2272 3819 2704
rect 3631 1409 3819 2272
rect 3889 3590 4077 4264
rect 3889 3169 3906 3590
rect 4059 3169 4077 3590
rect 3889 2194 4077 3169
rect 3889 1773 3906 2194
rect 4059 1773 4077 2194
rect 3373 -213 3390 208
rect 3543 -213 3561 208
rect 3373 -1188 3561 -213
rect 3373 -1609 3390 -1188
rect 3543 -1609 3561 -1188
rect 3373 -1741 3561 -1609
rect 3631 -686 3819 1241
rect 3631 -1107 3649 -686
rect 3802 -1107 3819 -686
rect 3631 -1741 3819 -1107
rect 3889 208 4077 1773
rect 4147 4100 4335 4264
rect 4147 3668 4162 4100
rect 4316 3668 4335 4100
rect 4147 2704 4335 3668
rect 4147 2272 4162 2704
rect 4316 2272 4335 2704
rect 4147 1409 4335 2272
rect 4405 3590 4593 4264
rect 4405 3169 4422 3590
rect 4575 3169 4593 3590
rect 4405 2194 4593 3169
rect 4405 1773 4422 2194
rect 4575 1773 4593 2194
rect 3889 -213 3906 208
rect 4059 -213 4077 208
rect 3889 -1188 4077 -213
rect 3889 -1609 3906 -1188
rect 4059 -1609 4077 -1188
rect 3889 -1741 4077 -1609
rect 4147 714 4335 1241
rect 4147 293 4165 714
rect 4318 293 4335 714
rect 4147 -1741 4335 293
rect 4405 208 4593 1773
rect 4405 -213 4422 208
rect 4575 -213 4593 208
rect 4405 -1188 4593 -213
rect 4405 -1609 4422 -1188
rect 4575 -1609 4593 -1188
rect 4405 -1741 4593 -1609
rect 4885 4229 4908 4324
rect 5291 4229 5314 4324
rect 4885 4099 5314 4229
rect 4885 3667 4898 4099
rect 5297 3667 5314 4099
rect 4885 2706 5314 3667
rect 4885 2279 4900 2706
rect 5295 2279 5314 2706
rect 4885 1609 5314 2279
rect 4885 1484 4898 1609
rect 5303 1484 5314 1609
rect 463 -3514 471 -3317
rect 636 -3514 650 -3317
rect 463 -3784 650 -3514
rect 4885 -2789 5314 1484
rect 4885 -2908 4901 -2789
rect 5299 -2908 5314 -2789
rect -305 -4309 -297 -4111
rect 112 -4309 124 -4111
rect -305 -4576 124 -4309
rect 4885 -4669 5314 -2908
rect 4885 -4805 4902 -4669
rect 5295 -4805 5314 -4669
rect 4885 -4821 5314 -4805
use pa_via  pa_via_0
timestamp 1718247345
transform 1 0 907 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_1
timestamp 1718247345
transform 1 0 138 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_2
timestamp 1718247345
transform 1 0 655 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_3
timestamp 1718247345
transform 1 0 1169 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_4
timestamp 1718247345
transform 1 0 395 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_5
timestamp 1718247345
transform 1 0 4346 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_6
timestamp 1718247345
transform 1 0 2023 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_7
timestamp 1718247345
transform 1 0 2282 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_8
timestamp 1718247345
transform 1 0 2542 0 1 -4717
box -10 3586 63 4043
use pa_via  pa_via_9
timestamp 1718247345
transform 1 0 2800 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_10
timestamp 1718247345
transform 1 0 3057 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_11
timestamp 1718247345
transform 1 0 3319 0 1 -5223
box -10 3586 63 4043
use pa_via  pa_via_12
timestamp 1718247345
transform 1 0 3574 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_13
timestamp 1718247345
transform 1 0 3831 0 1 -5222
box -10 3586 63 4043
use pa_via  pa_via_14
timestamp 1718247345
transform 1 0 4092 0 1 -4718
box -10 3586 63 4043
use pa_via  pa_via_15
timestamp 1718247345
transform 1 0 4608 0 1 -4717
box -10 3586 63 4043
use pa_via  pa_via_16
timestamp 1718247345
transform 1 0 902 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_17
timestamp 1718247345
transform 1 0 390 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_18
timestamp 1718247345
transform 1 0 1164 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_19
timestamp 1718247345
transform 1 0 650 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_20
timestamp 1718247345
transform 1 0 133 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_21
timestamp 1718247345
transform 1 0 3826 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_22
timestamp 1718247345
transform 1 0 3314 0 1 -435
box -10 3586 63 4043
use pa_via  pa_via_23
timestamp 1718247345
transform 1 0 2795 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_24
timestamp 1718247345
transform 1 0 2277 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_25
timestamp 1718247345
transform 1 0 4341 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_26
timestamp 1718247345
transform 1 0 4603 0 1 71
box -10 3586 63 4043
use pa_via  pa_via_27
timestamp 1718247345
transform 1 0 4087 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_28
timestamp 1718247345
transform 1 0 3569 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_29
timestamp 1718247345
transform 1 0 3052 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_30
timestamp 1718247345
transform 1 0 2537 0 1 71
box -10 3586 63 4043
use pa_via  pa_via_31
timestamp 1718247345
transform 1 0 2018 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_32
timestamp 1718247345
transform 1 0 135 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_33
timestamp 1718247345
transform 1 0 392 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_34
timestamp 1718247345
transform 1 0 652 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_35
timestamp 1718247345
transform 1 0 904 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_36
timestamp 1718247345
transform 1 0 1166 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_37
timestamp 1718247345
transform 1 0 2539 0 1 -1324
box -10 3586 63 4043
use pa_via  pa_via_38
timestamp 1718247345
transform 1 0 2797 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_39
timestamp 1718247345
transform 1 0 3054 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_40
timestamp 1718247345
transform 1 0 3316 0 1 -1830
box -10 3586 63 4043
use pa_via  pa_via_41
timestamp 1718247345
transform 1 0 3571 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_42
timestamp 1718247345
transform 1 0 3828 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_43
timestamp 1718247345
transform 1 0 4089 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_44
timestamp 1718247345
transform 1 0 4343 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_45
timestamp 1718247345
transform 1 0 4605 0 1 -1324
box -10 3586 63 4043
use pa_via  pa_via_46
timestamp 1718247345
transform 1 0 2020 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_47
timestamp 1718247345
transform 1 0 2279 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_48
timestamp 1718247345
transform 1 0 904 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_49
timestamp 1718247345
transform 1 0 392 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_50
timestamp 1718247345
transform 1 0 2279 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_51
timestamp 1718247345
transform 1 0 4343 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_52
timestamp 1718247345
transform 1 0 3828 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_53
timestamp 1718247345
transform 1 0 3316 0 1 -3817
box -10 3586 63 4043
use pa_via  pa_via_54
timestamp 1718247345
transform 1 0 2797 0 1 -3816
box -10 3586 63 4043
use pa_via  pa_via_55
timestamp 1718247345
transform 1 0 135 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_56
timestamp 1718247345
transform 1 0 1166 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_57
timestamp 1718247345
transform 1 0 652 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_58
timestamp 1718247345
transform 1 0 2020 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_59
timestamp 1718247345
transform 1 0 4605 0 1 -3311
box -10 3586 63 4043
use pa_via  pa_via_60
timestamp 1718247345
transform 1 0 4089 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_61
timestamp 1718247345
transform 1 0 3571 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_62
timestamp 1718247345
transform 1 0 3054 0 1 -3312
box -10 3586 63 4043
use pa_via  pa_via_63
timestamp 1718247345
transform 1 0 2539 0 1 -3311
box -10 3586 63 4043
use pa_via_short  pa_via_short_0
timestamp 1718247345
transform 1 0 -1878 0 1 -2428
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_1
timestamp 1718247345
transform 1 0 -3665 0 1 -1627
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_2
timestamp 1718247345
transform 0 1 4361 -1 0 2004
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_3
timestamp 1718247345
transform 1 0 -3510 0 1 -2175
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_4
timestamp 1718247345
transform 1 0 -2912 0 1 -2166
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_5
timestamp 1718247345
transform 1 0 -1718 0 1 -2168
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_6
timestamp 1718247345
transform 1 0 -1128 0 1 -2171
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_7
timestamp 1718247345
transform 1 0 -1291 0 1 -2426
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_8
timestamp 1718247345
transform 1 0 -3073 0 1 -1892
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_9
timestamp 1718247345
transform 0 1 4360 -1 0 2932
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_10
timestamp 1718247345
transform -1 0 6493 0 -1 -874
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_11
timestamp 1718247345
transform 0 1 3115 -1 0 6335
box 4944 -1889 5010 -1683
use sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y  sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y_0 paramcells
timestamp 1718247345
transform -1 0 3178 0 1 -3814
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  sky130_fd_pr__pfet_g5v0d10v5_FGL9FS_0 paramcells
timestamp 1718247345
transform -1 0 675 0 1 -1153
box -745 -797 745 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  sky130_fd_pr__pfet_g5v0d10v5_FGL9FS_1
timestamp 1718247345
transform -1 0 675 0 1 251
box -745 -797 745 797
use sky130_fd_sc_hvl__lsbuflv2hv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1718247345
transform -1 0 7769 0 1 -463
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  x2
timestamp 1718247345
transform -1 0 7769 0 1 1165
box -66 -43 2178 1671
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM1_1 paramcells
timestamp 1718247345
transform -1 0 3339 0 1 2245
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM1_2
timestamp 1718247345
transform -1 0 3339 0 1 3649
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  XM2_2
timestamp 1718247345
transform -1 0 675 0 1 3649
box -745 -797 745 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  XM3_2
timestamp 1718247345
transform -1 0 675 0 1 2245
box -745 -797 745 797
use sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y  XM4_2
timestamp 1718247345
transform -1 0 3770 0 1 -3814
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM5 paramcells
timestamp 1718247345
transform -1 0 1392 0 1 -3814
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM6_1
timestamp 1718247345
transform -1 0 3339 0 1 -1153
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM6_2
timestamp 1718247345
transform -1 0 3339 0 1 251
box -1519 -797 1519 797
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM8
timestamp 1718247345
transform -1 0 1986 0 1 -3814
box -278 -758 278 758
<< labels >>
flabel metal1 -280 2855 -80 3055 0 FreeSans 256 0 0 0 vinn
port 3 nsew
flabel metal1 -274 1237 -74 1437 0 FreeSans 256 0 0 0 vinp
port 4 nsew
flabel metal3 4973 4344 5173 4544 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal3 -230 -4547 -30 -4347 0 FreeSans 256 0 0 0 avss
port 7 nsew
flabel metal2 5116 -3705 5316 -3505 0 FreeSans 256 0 0 0 oneg
port 5 nsew
flabel metal2 5116 -3433 5316 -3233 0 FreeSans 256 0 0 0 opos
port 6 nsew
flabel metal2 7105 -566 7540 -477 0 FreeSans 800 0 0 0 dvss
port 9 nsew
flabel metal2 6471 -581 6906 -492 0 FreeSans 800 0 0 0 dvdd
port 8 nsew
flabel metal1 7642 1460 7842 1660 0 FreeSans 256 0 0 0 enab
port 1 nsew
flabel metal1 7630 -162 7830 38 0 FreeSans 256 0 0 0 clka
port 2 nsew
<< end >>
