** sch_path: /home/ttuser/chipalooza2024/sky130_icrg_ip__ulpcomp/cace/tb_voltage_swing.sch
**.subckt tb_voltage_swing
R1 vout net1 200k m=1
x1 dvdd avdd ena net2 net1 vout voutb avss dvss sky130_icrg_ip__ulpcomp
XC1 vout GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
V1 net2 avss 0.5 AC 0.9
avdd avdd GND DC {avdd}
dvdd dvdd GND DC {dvdd}
avss avss GND DC {avss}
dvss dvss GND DC {dvss}
ena ena GND Pulse(0 1.8 0 0.1n 0.1n 0.5n 1n)
**** begin user architecture code



.include {DUT_path}

.lib /home/ttuser/pdk/sky130A/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}

.option warn=1


.control
tran [1.0 / {frequency} / 100] [1 / {frequency}]
set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -V(vout)
quit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
