magic
tech sky130A
timestamp 1717166647
<< pwell >>
rect -139 -379 139 379
<< mvnmos >>
rect -25 -250 25 250
<< mvndiff >>
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
<< mvndiffc >>
rect -48 -244 -31 244
rect 31 -244 48 244
<< mvpsubdiff >>
rect -121 355 121 361
rect -121 338 -67 355
rect 67 338 121 355
rect -121 332 121 338
rect -121 307 -92 332
rect -121 -307 -115 307
rect -98 -307 -92 307
rect 92 307 121 332
rect -121 -332 -92 -307
rect 92 -307 98 307
rect 115 -307 121 307
rect 92 -332 121 -307
rect -121 -338 121 -332
rect -121 -355 -67 -338
rect 67 -355 121 -338
rect -121 -361 121 -355
<< mvpsubdiffcont >>
rect -67 338 67 355
rect -115 -307 -98 307
rect 98 -307 115 307
rect -67 -355 67 -338
<< poly >>
rect -25 286 25 294
rect -25 269 -17 286
rect 17 269 25 286
rect -25 250 25 269
rect -25 -269 25 -250
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -294 25 -286
<< polycont >>
rect -17 269 17 286
rect -17 -286 17 -269
<< locali >>
rect -115 338 -67 355
rect 67 338 115 355
rect -115 307 -98 338
rect 98 307 115 338
rect -25 269 -17 286
rect 17 269 25 286
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -115 -338 -98 -307
rect 98 -338 115 -307
rect -115 -355 -67 -338
rect 67 -355 115 -338
<< viali >>
rect -17 269 17 286
rect -48 -244 -31 244
rect 31 -244 48 244
rect -17 -286 17 -269
<< metal1 >>
rect -23 286 23 289
rect -23 269 -17 286
rect 17 269 23 286
rect -23 266 23 269
rect -51 244 -28 250
rect -51 -244 -48 244
rect -31 -244 -28 244
rect -51 -250 -28 -244
rect 28 244 51 250
rect 28 -244 31 244
rect 48 -244 51 244
rect 28 -250 51 -244
rect -23 -269 23 -266
rect -23 -286 -17 -269
rect 17 -286 23 -269
rect -23 -289 23 -286
<< properties >>
string FIXED_BBOX -106 -346 106 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
