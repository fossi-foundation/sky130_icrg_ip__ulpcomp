magic
tech sky130A
magscale 1 2
timestamp 1717166647
<< nwell >>
rect -487 -2415 487 2415
<< mvpmos >>
rect -229 118 -29 2118
rect 29 118 229 2118
rect -229 -2118 -29 -118
rect 29 -2118 229 -118
<< mvpdiff >>
rect -287 2106 -229 2118
rect -287 130 -275 2106
rect -241 130 -229 2106
rect -287 118 -229 130
rect -29 2106 29 2118
rect -29 130 -17 2106
rect 17 130 29 2106
rect -29 118 29 130
rect 229 2106 287 2118
rect 229 130 241 2106
rect 275 130 287 2106
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -2106 -275 -130
rect -241 -2106 -229 -130
rect -287 -2118 -229 -2106
rect -29 -130 29 -118
rect -29 -2106 -17 -130
rect 17 -2106 29 -130
rect -29 -2118 29 -2106
rect 229 -130 287 -118
rect 229 -2106 241 -130
rect 275 -2106 287 -130
rect 229 -2118 287 -2106
<< mvpdiffc >>
rect -275 130 -241 2106
rect -17 130 17 2106
rect 241 130 275 2106
rect -275 -2106 -241 -130
rect -17 -2106 17 -130
rect 241 -2106 275 -130
<< mvnsubdiff >>
rect -421 2337 421 2349
rect -421 2303 -313 2337
rect 313 2303 421 2337
rect -421 2291 421 2303
rect -421 2241 -363 2291
rect -421 -2241 -409 2241
rect -375 -2241 -363 2241
rect 363 2241 421 2291
rect -421 -2291 -363 -2241
rect 363 -2241 375 2241
rect 409 -2241 421 2241
rect 363 -2291 421 -2241
rect -421 -2303 421 -2291
rect -421 -2337 -313 -2303
rect 313 -2337 421 -2303
rect -421 -2349 421 -2337
<< mvnsubdiffcont >>
rect -313 2303 313 2337
rect -409 -2241 -375 2241
rect 375 -2241 409 2241
rect -313 -2337 313 -2303
<< poly >>
rect -229 2199 -29 2215
rect -229 2165 -213 2199
rect -45 2165 -29 2199
rect -229 2118 -29 2165
rect 29 2199 229 2215
rect 29 2165 45 2199
rect 213 2165 229 2199
rect 29 2118 229 2165
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -2165 -29 -2118
rect -229 -2199 -213 -2165
rect -45 -2199 -29 -2165
rect -229 -2215 -29 -2199
rect 29 -2165 229 -2118
rect 29 -2199 45 -2165
rect 213 -2199 229 -2165
rect 29 -2215 229 -2199
<< polycont >>
rect -213 2165 -45 2199
rect 45 2165 213 2199
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -2199 -45 -2165
rect 45 -2199 213 -2165
<< locali >>
rect -409 2303 -313 2337
rect 313 2303 409 2337
rect -409 2241 -375 2303
rect 375 2241 409 2303
rect -229 2165 -213 2199
rect -45 2165 -29 2199
rect 29 2165 45 2199
rect 213 2165 229 2199
rect -275 2106 -241 2122
rect -275 114 -241 130
rect -17 2106 17 2122
rect -17 114 17 130
rect 241 2106 275 2122
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -2122 -241 -2106
rect -17 -130 17 -114
rect -17 -2122 17 -2106
rect 241 -130 275 -114
rect 241 -2122 275 -2106
rect -229 -2199 -213 -2165
rect -45 -2199 -29 -2165
rect 29 -2199 45 -2165
rect 213 -2199 229 -2165
rect -409 -2303 -375 -2241
rect 375 -2303 409 -2241
rect -409 -2337 -313 -2303
rect 313 -2337 409 -2303
<< viali >>
rect -213 2165 -45 2199
rect 45 2165 213 2199
rect -275 130 -241 2106
rect -17 130 17 2106
rect 241 130 275 2106
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -2106 -241 -130
rect -17 -2106 17 -130
rect 241 -2106 275 -130
rect -213 -2199 -45 -2165
rect 45 -2199 213 -2165
<< metal1 >>
rect -225 2199 -33 2205
rect -225 2165 -213 2199
rect -45 2165 -33 2199
rect -225 2159 -33 2165
rect 33 2199 225 2205
rect 33 2165 45 2199
rect 213 2165 225 2199
rect 33 2159 225 2165
rect -281 2106 -235 2118
rect -281 130 -275 2106
rect -241 130 -235 2106
rect -281 118 -235 130
rect -23 2106 23 2118
rect -23 130 -17 2106
rect 17 130 23 2106
rect -23 118 23 130
rect 235 2106 281 2118
rect 235 130 241 2106
rect 275 130 281 2106
rect 235 118 281 130
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -130 -235 -118
rect -281 -2106 -275 -130
rect -241 -2106 -235 -130
rect -281 -2118 -235 -2106
rect -23 -130 23 -118
rect -23 -2106 -17 -130
rect 17 -2106 23 -130
rect -23 -2118 23 -2106
rect 235 -130 281 -118
rect 235 -2106 241 -130
rect 275 -2106 281 -130
rect 235 -2118 281 -2106
rect -225 -2165 -33 -2159
rect -225 -2199 -213 -2165
rect -45 -2199 -33 -2165
rect -225 -2205 -33 -2199
rect 33 -2165 225 -2159
rect 33 -2199 45 -2165
rect 213 -2199 225 -2165
rect 33 -2205 225 -2199
<< properties >>
string FIXED_BBOX -392 -2320 392 2320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
