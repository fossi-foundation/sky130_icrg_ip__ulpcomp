magic
tech sky130A
magscale 1 2
timestamp 1717203078
<< dnwell >>
rect 402 -4635 4688 -2706
<< nwell >>
rect 293 -2912 4797 -2583
rect 293 -4429 608 -2912
rect 2297 -4429 2865 -2912
rect 4482 -4429 4797 -2912
rect 293 -4744 4797 -4429
<< mvpsubdiff >>
rect 5434 2868 5494 2902
rect 7903 2868 7963 2902
rect 5434 2842 5468 2868
rect 5434 -534 5468 -508
rect 7929 2842 7963 2868
rect 7929 -534 7963 -508
rect 5434 -568 5494 -534
rect 7903 -568 7963 -534
<< mvnsubdiff >>
rect 359 -2689 4731 -2663
rect 359 -2710 456 -2689
rect 359 -4598 379 -2710
rect 413 -2725 456 -2710
rect 4616 -2725 4731 -2689
rect 413 -2737 4731 -2725
rect 413 -4598 433 -2737
rect 359 -4604 433 -4598
rect 4657 -2775 4731 -2737
rect 4657 -4598 4677 -2775
rect 4711 -4598 4731 -2775
rect 4657 -4604 4731 -4598
rect 359 -4624 4731 -4604
rect 359 -4658 439 -4624
rect 4651 -4658 4731 -4624
rect 359 -4678 4731 -4658
<< mvpsubdiffcont >>
rect 5494 2868 7903 2902
rect 5434 -508 5468 2842
rect 7929 -508 7963 2842
rect 5494 -568 7903 -534
<< mvnsubdiffcont >>
rect 379 -4598 413 -2710
rect 456 -2725 4616 -2689
rect 4677 -4598 4711 -2775
rect 439 -4658 4651 -4624
<< locali >>
rect 1797 4377 4706 4389
rect 1797 4340 1825 4377
rect 4634 4340 4706 4377
rect 1797 4317 4706 4340
rect 19 3148 160 4136
rect 1187 3146 1328 4134
rect 5434 2868 5494 2902
rect 7903 2868 7963 2902
rect 5434 2842 7963 2868
rect 22 1745 163 2733
rect 1190 1744 1331 2732
rect -6 1519 1347 1596
rect 1797 1560 4704 1583
rect 1797 1523 1833 1560
rect 4652 1523 4704 1560
rect 1797 1510 4704 1523
rect -3 1054 1350 1131
rect 1799 1118 4698 1128
rect 1799 1072 1826 1118
rect 4677 1072 4698 1118
rect 1799 1063 4698 1072
rect 21 -97 162 891
rect 1190 -92 1331 896
rect 5433 -508 5434 -455
rect 5468 2789 7929 2842
rect 5468 -455 5540 2789
rect 5640 2369 5745 2382
rect 5640 2162 5651 2369
rect 5732 2162 5745 2369
rect 5640 2149 5745 2162
rect 7270 1596 7472 1609
rect 7270 1490 7286 1596
rect 7458 1490 7472 1596
rect 7270 1475 7472 1490
rect 5641 738 5746 751
rect 5641 531 5652 738
rect 5733 531 5746 738
rect 5641 518 5746 531
rect 7270 -32 7472 -19
rect 7270 -138 7286 -32
rect 7458 -138 7472 -32
rect 7270 -153 7472 -138
rect 7858 -455 7929 2789
rect 5468 -508 7929 -455
rect 22 -1501 163 -513
rect 1188 -1501 1329 -513
rect 5433 -534 7963 -508
rect 5433 -563 5494 -534
rect 5434 -568 5494 -563
rect 7903 -568 7963 -534
rect -3 -1735 1350 -1658
rect 1792 -1673 4702 -1667
rect 1792 -1719 1826 -1673
rect 4677 -1719 4702 -1673
rect 1792 -1738 4702 -1719
rect 615 -2682 4711 -2667
rect 615 -2689 642 -2682
rect 379 -2710 456 -2689
rect 413 -2725 456 -2710
rect 4666 -2720 4711 -2682
rect 4616 -2725 4711 -2720
rect 615 -2736 4711 -2725
rect 4677 -2775 4711 -2736
rect 1119 -2947 2290 -2935
rect 1119 -2999 1153 -2947
rect 1119 -3019 2290 -2999
rect 1119 -3699 1178 -3019
rect 1119 -3708 1197 -3699
rect 1119 -3907 1133 -3708
rect 1185 -3907 1197 -3708
rect 1119 -3918 1197 -3907
rect 1119 -4313 1178 -3918
rect 1602 -4313 1772 -3019
rect 2201 -3702 2290 -3019
rect 2180 -3714 2290 -3702
rect 2180 -3907 2195 -3714
rect 2276 -3907 2290 -3714
rect 2180 -3917 2290 -3907
rect 2201 -4313 2290 -3917
rect 1119 -4329 2290 -4313
rect 1119 -4381 1163 -4329
rect 1119 -4397 2290 -4381
rect 2855 -2947 4041 -2935
rect 4009 -2999 4041 -2947
rect 2855 -3019 4041 -2999
rect 2855 -3968 2971 -3019
rect 2855 -4161 2867 -3968
rect 2968 -4161 2971 -3968
rect 2855 -4313 2971 -4161
rect 3394 -4313 3564 -3019
rect 3982 -4313 4041 -3019
rect 2855 -4329 4041 -4313
rect 4019 -4381 4041 -4329
rect 2855 -4397 4041 -4381
rect 379 -4602 413 -4598
rect 4677 -4602 4711 -4598
rect 371 -4619 4720 -4602
rect 371 -4660 388 -4619
rect 4681 -4660 4720 -4619
rect 371 -4677 4720 -4660
<< viali >>
rect 1825 4340 4634 4377
rect 1833 1523 4652 1560
rect 1826 1072 4677 1118
rect 5651 2162 5732 2369
rect 7286 1490 7458 1596
rect 5652 531 5733 738
rect 7286 -138 7458 -32
rect 1826 -1719 4677 -1673
rect 642 -2689 4666 -2682
rect 642 -2720 4616 -2689
rect 4616 -2720 4666 -2689
rect 1153 -2999 2290 -2947
rect 1133 -3907 1185 -3708
rect 2195 -3907 2276 -3714
rect 1163 -4381 2290 -4329
rect 2855 -2999 4009 -2947
rect 2867 -4161 2968 -3968
rect 2855 -4381 4019 -4329
rect 388 -4624 4681 -4619
rect 388 -4658 439 -4624
rect 439 -4658 4651 -4624
rect 4651 -4658 4681 -4624
rect 388 -4660 4681 -4658
<< metal1 >>
rect 1797 4377 5224 4388
rect 1797 4340 1825 4377
rect 4634 4340 5224 4377
rect 1797 4324 5224 4340
rect 1797 4317 4818 4324
rect 4795 4229 4818 4317
rect 5201 4229 5224 4324
rect -280 2971 -80 3055
rect 275 2971 322 4226
rect 533 2971 580 4226
rect 791 2971 838 4226
rect 1049 2971 1096 4226
rect -280 2923 1546 2971
rect 2067 2961 2114 4223
rect 2325 2961 2372 4223
rect 2583 2961 2630 4223
rect 2841 2961 2888 4223
rect 3099 2961 3146 4223
rect 3357 2961 3404 4223
rect 3615 2961 3662 4223
rect 3873 2961 3920 4223
rect 4131 2961 4178 4223
rect 4389 2961 4436 4223
rect 4795 4211 5224 4229
rect -280 2922 248 2923
rect -280 2855 -80 2922
rect 275 1733 322 2832
rect 533 1751 580 2832
rect 791 1786 838 2832
rect 271 1681 322 1733
rect 529 1681 580 1751
rect 787 1681 838 1786
rect 1049 1746 1096 2832
rect 1045 1681 1096 1746
rect -274 1380 -74 1437
rect 271 1380 318 1681
rect 529 1380 576 1681
rect 787 1380 834 1681
rect 1045 1380 1092 1681
rect -274 1332 1397 1380
rect -274 1237 -74 1332
rect 1484 1275 1546 2923
rect 2062 2919 4896 2961
rect 2067 1678 2114 2919
rect 2325 1678 2372 2919
rect 2583 1678 2630 2919
rect 2841 1678 2888 2919
rect 3099 1678 3146 2919
rect 3357 1678 3404 2919
rect 3615 1678 3662 2919
rect 3873 1678 3920 2919
rect 4131 1678 4178 2919
rect 4389 1678 4436 2919
rect 4854 2255 4896 2919
rect 5450 2799 7948 2903
rect 5450 2691 7130 2799
rect 7520 2691 7948 2799
rect 5450 2672 7948 2691
rect 5640 2369 5745 2382
rect 5640 2255 5651 2369
rect 4854 2210 5651 2255
rect 4896 2207 5651 2210
rect 5640 2162 5651 2207
rect 5732 2162 5745 2369
rect 5640 2149 5745 2162
rect 5661 1894 5867 2064
rect 6261 1894 7765 2064
rect 4795 1609 5224 1619
rect 4795 1581 4808 1609
rect 1797 1560 4808 1581
rect 1797 1523 1833 1560
rect 4652 1523 4808 1560
rect 1797 1510 4808 1523
rect 4795 1484 4808 1510
rect 5213 1484 5224 1609
rect 4795 1473 5224 1484
rect 7270 1596 7472 1609
rect 7270 1490 7286 1596
rect 7458 1573 7472 1596
rect 7642 1573 7842 1664
rect 7458 1517 7842 1573
rect 7458 1490 7472 1517
rect 7270 1475 7472 1490
rect 7642 1464 7842 1517
rect 271 1227 1546 1275
rect 271 -182 318 1227
rect 529 -182 576 1227
rect 787 -182 834 1227
rect 1045 -182 1092 1227
rect 1796 1118 4744 1149
rect 1484 -289 1546 1103
rect 1796 1072 1826 1118
rect 4677 1072 4744 1118
rect 5653 1080 7137 1250
rect 7511 1080 7757 1250
rect 1796 1048 4744 1072
rect 2063 -286 2110 959
rect 2321 -286 2368 959
rect 2579 -286 2626 959
rect 2837 -286 2884 959
rect 3095 -286 3142 959
rect 3353 -286 3400 959
rect 3611 -286 3658 959
rect 3869 -286 3916 959
rect 4127 -286 4174 959
rect 4385 -286 4432 959
rect 4652 366 4744 1048
rect 5641 738 5746 751
rect 5641 657 5652 738
rect 4652 -71 4664 366
rect 4736 -71 4744 366
rect 4652 -81 4744 -71
rect 5294 609 5652 657
rect 5294 -216 5336 609
rect 5641 531 5652 609
rect 5733 531 5746 738
rect 5641 518 5746 531
rect 5659 262 5866 432
rect 6260 262 7763 432
rect 7270 -32 7472 -19
rect 7270 -138 7286 -32
rect 7458 -51 7472 -32
rect 7630 -51 7830 42
rect 7458 -107 7830 -51
rect 7458 -138 7472 -107
rect 7270 -153 7472 -138
rect 7630 -158 7830 -107
rect 5294 -286 5334 -216
rect 249 -322 1546 -289
rect 271 -1583 318 -322
rect 529 -1583 576 -322
rect 787 -1583 834 -322
rect 1045 -1583 1092 -322
rect 2056 -328 5334 -286
rect 2063 -1586 2110 -328
rect 2321 -1586 2368 -328
rect 2579 -1586 2626 -328
rect 2837 -1586 2884 -328
rect 3095 -1586 3142 -328
rect 3353 -1586 3400 -328
rect 3611 -1586 3658 -328
rect 3869 -1586 3916 -328
rect 4127 -1586 4174 -328
rect 4385 -1586 4432 -328
rect 4649 -1040 4748 -1025
rect 4649 -1483 4657 -1040
rect 4739 -1483 4748 -1040
rect 4649 -1658 4748 -1483
rect 1780 -1673 4748 -1658
rect 1780 -1719 1826 -1673
rect 4677 -1719 4748 -1673
rect 1780 -1759 4748 -1719
rect 5294 -1878 5334 -328
rect 5653 -467 7121 -366
rect 7519 -467 7765 -366
rect 5653 -470 7765 -467
rect 2640 -1918 5334 -1878
rect 4795 -2645 5224 -2634
rect 4795 -2669 4811 -2645
rect 615 -2682 4811 -2669
rect 615 -2720 642 -2682
rect 4666 -2720 4811 -2682
rect 615 -2736 4811 -2720
rect 4795 -2764 4811 -2736
rect 5209 -2764 5224 -2645
rect 4795 -2776 5224 -2764
rect 1121 -2947 2315 -2932
rect 1121 -2999 1153 -2947
rect 2290 -2999 2315 -2947
rect 1121 -3021 2315 -2999
rect 2550 -3068 2596 -2803
rect 2828 -2947 4040 -2932
rect 2828 -2999 2855 -2947
rect 4009 -2999 4040 -2947
rect 2828 -3012 2871 -2999
rect 3953 -3012 4040 -2999
rect 2828 -3021 4040 -3012
rect 1344 -3109 2596 -3068
rect 3128 -3109 3872 -3068
rect 1120 -3708 1197 -3699
rect 1120 -3907 1133 -3708
rect 1185 -3907 1197 -3708
rect 1120 -3918 1197 -3907
rect 1371 -4233 1408 -3112
rect 1965 -4235 2002 -3114
rect 3195 -3116 3280 -3109
rect 3787 -3114 3872 -3109
rect 3158 -3138 3280 -3116
rect 2180 -3714 2289 -3702
rect 2180 -3907 2195 -3714
rect 2276 -3907 2289 -3714
rect 2180 -3917 2289 -3907
rect 2855 -3968 2982 -3958
rect 2855 -4161 2867 -3968
rect 2968 -4161 2982 -3968
rect 2855 -4174 2982 -4161
rect 3158 -4237 3195 -3138
rect 3234 -3187 3280 -3138
rect 3752 -3138 3872 -3114
rect 3752 -4235 3789 -3138
rect 3826 -3177 3872 -3138
rect 1121 -4329 2315 -4313
rect 1121 -4381 1163 -4329
rect 2290 -4381 2315 -4329
rect 1121 -4397 2315 -4381
rect 2828 -4329 4043 -4313
rect 2828 -4381 2855 -4329
rect 4019 -4381 4043 -4329
rect 2828 -4397 4043 -4381
rect 4795 -4525 5224 -4509
rect 4795 -4602 4812 -4525
rect 371 -4619 4812 -4602
rect 371 -4660 388 -4619
rect 4681 -4660 4812 -4619
rect 371 -4661 4812 -4660
rect 5205 -4661 5224 -4525
rect 371 -4677 5224 -4661
<< via1 >>
rect 4818 4229 5201 4324
rect 7130 2691 7520 2799
rect 5867 1875 6261 2091
rect 6494 1773 6882 1830
rect 4808 1484 5213 1609
rect 7137 1076 7511 1261
rect 4664 -71 4736 366
rect 5866 248 6260 464
rect 6494 145 6882 202
rect 4657 -1483 4739 -1040
rect 7121 -467 7519 -356
rect 4811 -2764 5209 -2645
rect 2871 -2999 3953 -2947
rect 2871 -3012 3953 -2999
rect 1133 -3907 1185 -3708
rect 2195 -3907 2276 -3714
rect 2867 -4161 2968 -3968
rect 4812 -4661 5205 -4525
<< metal2 >>
rect 4795 4324 5224 4342
rect 4795 4229 4818 4324
rect 5201 4229 5224 4324
rect 4795 4211 5224 4229
rect 116 4106 1728 4115
rect 116 3674 982 4106
rect 1140 3674 1728 4106
rect 116 3656 1728 3674
rect 1928 4100 5225 4115
rect 1928 3668 2008 4100
rect 2162 3668 2524 4100
rect 2678 3668 3040 4100
rect 3194 3668 3556 4100
rect 3710 3668 4072 4100
rect 4226 4099 5225 4100
rect 4226 3668 4808 4099
rect 1928 3667 4808 3668
rect 5207 3667 5225 4099
rect 1928 3656 5225 3667
rect 116 3596 1726 3610
rect 116 3164 478 3596
rect 636 3164 1726 3596
rect 116 3151 1726 3164
rect 1921 3590 4590 3610
rect 1921 3169 2268 3590
rect 2421 3169 2784 3590
rect 2937 3169 3300 3590
rect 3453 3169 3816 3590
rect 3969 3169 4332 3590
rect 4485 3169 4590 3590
rect 1921 3151 4590 3169
rect 116 2719 1726 2722
rect 116 2287 729 2719
rect 887 2718 1726 2719
rect 1928 2721 5375 2722
rect 5849 2721 6284 2873
rect 887 2287 1728 2718
rect 116 2263 1728 2287
rect 1925 2261 1927 2718
rect 1928 2706 6284 2721
rect 1928 2704 4810 2706
rect 1928 2272 2008 2704
rect 2162 2272 2524 2704
rect 2678 2272 3040 2704
rect 3194 2272 3556 2704
rect 3710 2272 4072 2704
rect 4226 2279 4810 2704
rect 5205 2279 6284 2706
rect 4226 2272 6284 2279
rect 1928 2263 6284 2272
rect 4578 2262 6284 2263
rect 116 2209 1726 2215
rect 116 1777 224 2209
rect 382 1777 1726 2209
rect 1925 2194 4590 2215
rect 1925 2179 2268 2194
rect 116 1756 1726 1777
rect 1921 1773 2268 2179
rect 2421 1773 2784 2194
rect 2937 1773 3300 2194
rect 3453 1773 3816 2194
rect 3969 1773 4332 2194
rect 4485 1773 4590 2194
rect 1921 1756 4590 1773
rect 5849 2091 6284 2262
rect 5849 1875 5867 2091
rect 6261 1875 6284 2091
rect 4795 1609 5224 1619
rect 4795 1484 4808 1609
rect 5213 1484 5224 1609
rect 4795 1473 5224 1484
rect 1418 1325 1549 1391
rect 1482 1144 1549 1325
rect 1485 1143 1547 1144
rect 116 866 4597 879
rect 116 434 979 866
rect 1137 863 4597 866
rect 1137 442 2011 863
rect 2164 442 3045 863
rect 3198 860 4597 863
rect 3198 442 4075 860
rect 1137 439 4075 442
rect 4228 439 4597 860
rect 1137 434 4597 439
rect 116 420 4597 434
rect 5849 464 6284 1875
rect 116 367 1728 375
rect 116 -65 474 367
rect 632 -65 1728 367
rect 116 -84 1728 -65
rect 1928 366 4745 375
rect 1928 354 4664 366
rect 1928 -67 2268 354
rect 2421 -67 2784 354
rect 2937 -67 3300 354
rect 3453 -67 3816 354
rect 3969 -67 4332 354
rect 4485 -67 4664 354
rect 1928 -71 4664 -67
rect 4736 -71 4745 366
rect 1928 -84 4745 -71
rect 5849 248 5866 464
rect 6260 248 6284 464
rect 116 -540 4590 -527
rect 116 -542 3559 -540
rect 116 -974 728 -542
rect 886 -552 3559 -542
rect 886 -973 2525 -552
rect 2678 -961 3559 -552
rect 3712 -961 4590 -540
rect 5849 -577 6284 248
rect 6471 1830 6906 2874
rect 6471 1773 6494 1830
rect 6882 1773 6906 1830
rect 6471 202 6906 1773
rect 6471 145 6494 202
rect 6882 145 6906 202
rect 6471 -592 6906 145
rect 7105 2799 7540 2857
rect 7105 2691 7130 2799
rect 7520 2691 7540 2799
rect 7105 1261 7540 2691
rect 7105 1076 7137 1261
rect 7511 1076 7540 1261
rect 7105 -356 7540 1076
rect 7105 -467 7121 -356
rect 7519 -467 7540 -356
rect 7105 -562 7540 -467
rect 2678 -973 4590 -961
rect 886 -974 4590 -973
rect 116 -986 4590 -974
rect 116 -1044 1728 -1031
rect 116 -1476 227 -1044
rect 385 -1476 1728 -1044
rect 116 -1490 1728 -1476
rect 1928 -1040 4750 -1031
rect 1928 -1042 4657 -1040
rect 1928 -1463 2268 -1042
rect 2421 -1463 2784 -1042
rect 2937 -1463 3300 -1042
rect 3453 -1463 3816 -1042
rect 3969 -1463 4332 -1042
rect 4485 -1463 4657 -1042
rect 1928 -1483 4657 -1463
rect 4739 -1483 4750 -1040
rect 1928 -1490 4750 -1483
rect 2541 -2824 2598 -1916
rect 4795 -2645 5224 -2634
rect 4795 -2764 4811 -2645
rect 5209 -2764 5224 -2645
rect 4795 -2776 5224 -2764
rect -303 -2943 4049 -2931
rect -303 -3089 -283 -2943
rect 105 -2947 4049 -2943
rect 105 -3012 2871 -2947
rect 3953 -3012 4049 -2947
rect 105 -3089 4049 -3012
rect -303 -3109 4049 -3089
rect 210 -3173 3892 -3164
rect 210 -3370 471 -3173
rect 636 -3278 3892 -3173
rect 5026 -3278 5226 -3233
rect 636 -3370 5226 -3278
rect 210 -3374 5226 -3370
rect 210 -3379 3892 -3374
rect 210 -3437 3897 -3426
rect 5026 -3433 5226 -3374
rect 210 -3634 221 -3437
rect 386 -3505 3897 -3437
rect 386 -3601 5226 -3505
rect 386 -3634 3897 -3601
rect 210 -3641 3897 -3634
rect 1102 -3708 3893 -3702
rect 5026 -3705 5226 -3601
rect 1102 -3907 1133 -3708
rect 1185 -3714 3893 -3708
rect 1185 -3907 2195 -3714
rect 2276 -3907 3893 -3714
rect 1102 -3918 3893 -3907
rect -305 -3967 3888 -3958
rect -305 -4165 -297 -3967
rect 112 -3968 3888 -3967
rect 112 -4161 2867 -3968
rect 2968 -4161 3888 -3968
rect 112 -4165 3888 -4161
rect -305 -4174 3888 -4165
rect 4795 -4525 5224 -4509
rect 4795 -4661 4812 -4525
rect 5205 -4661 5224 -4525
rect 4795 -4677 5224 -4661
<< via2 >>
rect 4818 4229 5201 4324
rect 982 3674 1140 4106
rect 2008 3668 2162 4100
rect 2524 3668 2678 4100
rect 3040 3668 3194 4100
rect 3556 3668 3710 4100
rect 4072 3668 4226 4100
rect 4808 3667 5207 4099
rect 478 3164 636 3596
rect 2268 3169 2421 3590
rect 2784 3169 2937 3590
rect 3300 3169 3453 3590
rect 3816 3169 3969 3590
rect 4332 3169 4485 3590
rect 729 2287 887 2719
rect 2008 2272 2162 2704
rect 2524 2272 2678 2704
rect 3040 2272 3194 2704
rect 3556 2272 3710 2704
rect 4072 2272 4226 2704
rect 4810 2279 5205 2706
rect 224 1777 382 2209
rect 2268 1773 2421 2194
rect 2784 1773 2937 2194
rect 3300 1773 3453 2194
rect 3816 1773 3969 2194
rect 4332 1773 4485 2194
rect 4808 1484 5213 1609
rect 979 434 1137 866
rect 2011 442 2164 863
rect 3045 442 3198 863
rect 4075 439 4228 860
rect 474 -65 632 367
rect 2268 -67 2421 354
rect 2784 -67 2937 354
rect 3300 -67 3453 354
rect 3816 -67 3969 354
rect 4332 -67 4485 354
rect 728 -974 886 -542
rect 2525 -973 2678 -552
rect 3559 -961 3712 -540
rect 227 -1476 385 -1044
rect 2268 -1463 2421 -1042
rect 2784 -1463 2937 -1042
rect 3300 -1463 3453 -1042
rect 3816 -1463 3969 -1042
rect 4332 -1463 4485 -1042
rect 4811 -2764 5209 -2645
rect -283 -3089 105 -2943
rect 471 -3370 636 -3173
rect 221 -3634 386 -3437
rect -297 -4165 112 -3967
rect 4812 -4661 5205 -4525
<< metal3 >>
rect -305 -2931 124 4434
rect 4795 4324 5224 4550
rect 211 2209 398 4262
rect 211 1777 224 2209
rect 382 1777 398 2209
rect 211 -1044 398 1777
rect 211 -1476 227 -1044
rect 385 -1476 398 -1044
rect -305 -2943 125 -2931
rect -305 -3089 -283 -2943
rect 105 -3089 125 -2943
rect -305 -3109 125 -3089
rect -305 -3967 124 -3109
rect 211 -3437 398 -1476
rect 211 -3634 221 -3437
rect 386 -3634 398 -3437
rect 211 -3642 398 -3634
rect 463 3596 650 4262
rect 463 3164 478 3596
rect 636 3164 650 3596
rect 463 367 650 3164
rect 463 -65 474 367
rect 632 -65 650 367
rect 463 -3173 650 -65
rect 715 2719 902 4262
rect 715 2287 729 2719
rect 887 2287 902 2719
rect 715 -542 902 2287
rect 715 -974 728 -542
rect 886 -974 902 -542
rect 715 -1615 902 -974
rect 967 4106 1154 4262
rect 967 3674 982 4106
rect 1140 3674 1154 4106
rect 967 866 1154 3674
rect 1993 4100 2181 4264
rect 1993 3668 2008 4100
rect 2162 3668 2181 4100
rect 1993 2704 2181 3668
rect 1993 2272 2008 2704
rect 2162 2272 2181 2704
rect 1993 1409 2181 2272
rect 2251 3590 2439 4264
rect 2251 3169 2268 3590
rect 2421 3169 2439 3590
rect 2251 2194 2439 3169
rect 2251 1773 2268 2194
rect 2421 1773 2439 2194
rect 967 434 979 866
rect 1137 434 1154 866
rect 967 -1615 1154 434
rect 1993 863 2181 1241
rect 1993 442 2011 863
rect 2164 442 2181 863
rect 1993 -1595 2181 442
rect 2251 354 2439 1773
rect 2509 4100 2697 4264
rect 2509 3668 2524 4100
rect 2678 3668 2697 4100
rect 2509 2704 2697 3668
rect 2509 2272 2524 2704
rect 2678 2272 2697 2704
rect 2509 1409 2697 2272
rect 2767 3590 2955 4264
rect 2767 3169 2784 3590
rect 2937 3169 2955 3590
rect 2767 2194 2955 3169
rect 2767 1773 2784 2194
rect 2937 1773 2955 2194
rect 2251 -67 2268 354
rect 2421 -67 2439 354
rect 2251 -1042 2439 -67
rect 2251 -1463 2268 -1042
rect 2421 -1463 2439 -1042
rect 2251 -1595 2439 -1463
rect 2509 -552 2697 1241
rect 2509 -973 2525 -552
rect 2678 -973 2697 -552
rect 2509 -1595 2697 -973
rect 2767 354 2955 1773
rect 3025 4100 3213 4264
rect 3025 3668 3040 4100
rect 3194 3668 3213 4100
rect 3025 2704 3213 3668
rect 3025 2272 3040 2704
rect 3194 2272 3213 2704
rect 3025 1409 3213 2272
rect 3283 3590 3471 4264
rect 3283 3169 3300 3590
rect 3453 3169 3471 3590
rect 3283 2194 3471 3169
rect 3283 1773 3300 2194
rect 3453 1773 3471 2194
rect 2767 -67 2784 354
rect 2937 -67 2955 354
rect 2767 -1042 2955 -67
rect 2767 -1463 2784 -1042
rect 2937 -1463 2955 -1042
rect 2767 -1595 2955 -1463
rect 3025 863 3213 1241
rect 3025 442 3045 863
rect 3198 442 3213 863
rect 3025 -1595 3213 442
rect 3283 354 3471 1773
rect 3541 4100 3729 4264
rect 3541 3668 3556 4100
rect 3710 3668 3729 4100
rect 3541 2704 3729 3668
rect 3541 2272 3556 2704
rect 3710 2272 3729 2704
rect 3541 1409 3729 2272
rect 3799 3590 3987 4264
rect 3799 3169 3816 3590
rect 3969 3169 3987 3590
rect 3799 2194 3987 3169
rect 3799 1773 3816 2194
rect 3969 1773 3987 2194
rect 3283 -67 3300 354
rect 3453 -67 3471 354
rect 3283 -1042 3471 -67
rect 3283 -1463 3300 -1042
rect 3453 -1463 3471 -1042
rect 3283 -1595 3471 -1463
rect 3541 -540 3729 1241
rect 3541 -961 3559 -540
rect 3712 -961 3729 -540
rect 3541 -1595 3729 -961
rect 3799 354 3987 1773
rect 4057 4100 4245 4264
rect 4057 3668 4072 4100
rect 4226 3668 4245 4100
rect 4057 2704 4245 3668
rect 4057 2272 4072 2704
rect 4226 2272 4245 2704
rect 4057 1409 4245 2272
rect 4315 3590 4503 4264
rect 4315 3169 4332 3590
rect 4485 3169 4503 3590
rect 4315 2194 4503 3169
rect 4315 1773 4332 2194
rect 4485 1773 4503 2194
rect 3799 -67 3816 354
rect 3969 -67 3987 354
rect 3799 -1042 3987 -67
rect 3799 -1463 3816 -1042
rect 3969 -1463 3987 -1042
rect 3799 -1595 3987 -1463
rect 4057 860 4245 1241
rect 4057 439 4075 860
rect 4228 439 4245 860
rect 4057 -1595 4245 439
rect 4315 354 4503 1773
rect 4315 -67 4332 354
rect 4485 -67 4503 354
rect 4315 -1042 4503 -67
rect 4315 -1463 4332 -1042
rect 4485 -1463 4503 -1042
rect 4315 -1595 4503 -1463
rect 4795 4229 4818 4324
rect 5201 4229 5224 4324
rect 4795 4099 5224 4229
rect 4795 3667 4808 4099
rect 5207 3667 5224 4099
rect 4795 2706 5224 3667
rect 4795 2279 4810 2706
rect 5205 2279 5224 2706
rect 4795 1609 5224 2279
rect 4795 1484 4808 1609
rect 5213 1484 5224 1609
rect 463 -3370 471 -3173
rect 636 -3370 650 -3173
rect 463 -3640 650 -3370
rect 4795 -2645 5224 1484
rect 4795 -2764 4811 -2645
rect 5209 -2764 5224 -2645
rect -305 -4165 -297 -3967
rect 112 -4165 124 -3967
rect -305 -4432 124 -4165
rect 4795 -4525 5224 -2764
rect 4795 -4661 4812 -4525
rect 5205 -4661 5224 -4525
rect 4795 -4677 5224 -4661
use pa_via  pa_via_0
timestamp 1717165164
transform 1 0 907 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_1
timestamp 1717165164
transform 1 0 138 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_2
timestamp 1717165164
transform 1 0 655 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_3
timestamp 1717165164
transform 1 0 1169 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_4
timestamp 1717165164
transform 1 0 395 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_5
timestamp 1717165164
transform 1 0 4256 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_6
timestamp 1717165164
transform 1 0 1933 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_7
timestamp 1717165164
transform 1 0 2192 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_8
timestamp 1717165164
transform 1 0 2452 0 1 -4571
box -10 3586 63 4043
use pa_via  pa_via_9
timestamp 1717165164
transform 1 0 2710 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_10
timestamp 1717165164
transform 1 0 2967 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_11
timestamp 1717165164
transform 1 0 3229 0 1 -5077
box -10 3586 63 4043
use pa_via  pa_via_12
timestamp 1717165164
transform 1 0 3484 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_13
timestamp 1717165164
transform 1 0 3741 0 1 -5076
box -10 3586 63 4043
use pa_via  pa_via_14
timestamp 1717165164
transform 1 0 4002 0 1 -4572
box -10 3586 63 4043
use pa_via  pa_via_15
timestamp 1717165164
transform 1 0 4518 0 1 -4571
box -10 3586 63 4043
use pa_via  pa_via_16
timestamp 1717165164
transform 1 0 902 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_17
timestamp 1717165164
transform 1 0 390 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_18
timestamp 1717165164
transform 1 0 1164 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_19
timestamp 1717165164
transform 1 0 650 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_20
timestamp 1717165164
transform 1 0 133 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_21
timestamp 1717165164
transform 1 0 3736 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_22
timestamp 1717165164
transform 1 0 3224 0 1 -435
box -10 3586 63 4043
use pa_via  pa_via_23
timestamp 1717165164
transform 1 0 2705 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_24
timestamp 1717165164
transform 1 0 2187 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_25
timestamp 1717165164
transform 1 0 4251 0 1 -434
box -10 3586 63 4043
use pa_via  pa_via_26
timestamp 1717165164
transform 1 0 4513 0 1 71
box -10 3586 63 4043
use pa_via  pa_via_27
timestamp 1717165164
transform 1 0 3997 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_28
timestamp 1717165164
transform 1 0 3479 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_29
timestamp 1717165164
transform 1 0 2962 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_30
timestamp 1717165164
transform 1 0 2447 0 1 71
box -10 3586 63 4043
use pa_via  pa_via_31
timestamp 1717165164
transform 1 0 1928 0 1 70
box -10 3586 63 4043
use pa_via  pa_via_32
timestamp 1717165164
transform 1 0 135 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_33
timestamp 1717165164
transform 1 0 392 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_34
timestamp 1717165164
transform 1 0 652 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_35
timestamp 1717165164
transform 1 0 904 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_36
timestamp 1717165164
transform 1 0 1166 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_37
timestamp 1717165164
transform 1 0 2449 0 1 -1324
box -10 3586 63 4043
use pa_via  pa_via_38
timestamp 1717165164
transform 1 0 2707 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_39
timestamp 1717165164
transform 1 0 2964 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_40
timestamp 1717165164
transform 1 0 3226 0 1 -1830
box -10 3586 63 4043
use pa_via  pa_via_41
timestamp 1717165164
transform 1 0 3481 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_42
timestamp 1717165164
transform 1 0 3738 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_43
timestamp 1717165164
transform 1 0 3999 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_44
timestamp 1717165164
transform 1 0 4253 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_45
timestamp 1717165164
transform 1 0 4515 0 1 -1324
box -10 3586 63 4043
use pa_via  pa_via_46
timestamp 1717165164
transform 1 0 1930 0 1 -1325
box -10 3586 63 4043
use pa_via  pa_via_47
timestamp 1717165164
transform 1 0 2189 0 1 -1829
box -10 3586 63 4043
use pa_via  pa_via_48
timestamp 1717165164
transform 1 0 904 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_49
timestamp 1717165164
transform 1 0 392 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_50
timestamp 1717165164
transform 1 0 2189 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_51
timestamp 1717165164
transform 1 0 4253 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_52
timestamp 1717165164
transform 1 0 3738 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_53
timestamp 1717165164
transform 1 0 3226 0 1 -3671
box -10 3586 63 4043
use pa_via  pa_via_54
timestamp 1717165164
transform 1 0 2707 0 1 -3670
box -10 3586 63 4043
use pa_via  pa_via_55
timestamp 1717165164
transform 1 0 135 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_56
timestamp 1717165164
transform 1 0 1166 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_57
timestamp 1717165164
transform 1 0 652 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_58
timestamp 1717165164
transform 1 0 1930 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_59
timestamp 1717165164
transform 1 0 4515 0 1 -3165
box -10 3586 63 4043
use pa_via  pa_via_60
timestamp 1717165164
transform 1 0 3999 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_61
timestamp 1717165164
transform 1 0 3481 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_62
timestamp 1717165164
transform 1 0 2964 0 1 -3166
box -10 3586 63 4043
use pa_via  pa_via_63
timestamp 1717165164
transform 1 0 2449 0 1 -3165
box -10 3586 63 4043
use pa_via_short  pa_via_short_0
timestamp 1717168741
transform 1 0 -1878 0 1 -2284
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_1
timestamp 1717168741
transform 1 0 -3665 0 1 -1483
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_2
timestamp 1717168741
transform 0 1 4361 -1 0 2148
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_3
timestamp 1717168741
transform 1 0 -3510 0 1 -2031
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_4
timestamp 1717168741
transform 1 0 -2912 0 1 -2022
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_5
timestamp 1717168741
transform 1 0 -1718 0 1 -2024
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_6
timestamp 1717168741
transform 1 0 -1128 0 1 -2027
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_7
timestamp 1717168741
transform 1 0 -1291 0 1 -2282
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_8
timestamp 1717168741
transform 1 0 -3073 0 1 -1748
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_9
timestamp 1717168741
transform 0 1 4360 -1 0 3078
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_10
timestamp 1717168741
transform -1 0 6493 0 -1 -728
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_11
timestamp 1717168741
transform 0 1 3115 -1 0 6335
box 4944 -1889 5010 -1683
use sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y  sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y_0 paramcells
timestamp 1717166647
transform -1 0 3178 0 1 -3670
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  sky130_fd_pr__pfet_g5v0d10v5_FGL9FS_0 paramcells
timestamp 1717166647
transform -1 0 675 0 1 -1007
box -745 -797 745 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  sky130_fd_pr__pfet_g5v0d10v5_FGL9FS_1
timestamp 1717166647
transform -1 0 675 0 1 397
box -745 -797 745 797
use sky130_fd_sc_hvl__lsbuflv2hv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform -1 0 7769 0 1 -459
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  x2
timestamp 1715205430
transform -1 0 7769 0 1 1169
box -66 -43 2178 1671
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM1_1 paramcells
timestamp 1717166647
transform -1 0 3249 0 1 2245
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM1_2
timestamp 1717166647
transform -1 0 3249 0 1 3649
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  XM2_2
timestamp 1717166647
transform -1 0 675 0 1 3649
box -745 -797 745 797
use sky130_fd_pr__pfet_g5v0d10v5_FGL9FS  XM3_2
timestamp 1717166647
transform -1 0 675 0 1 2245
box -745 -797 745 797
use sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y  XM4_2
timestamp 1717166647
transform -1 0 3770 0 1 -3670
box -278 -758 278 758
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM5 paramcells
timestamp 1717166647
transform -1 0 1392 0 1 -3670
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM6_1
timestamp 1717166647
transform -1 0 3249 0 1 -1007
box -1519 -797 1519 797
use sky130_fd_pr__pfet_g5v0d10v5_E2TVSU  XM6_2
timestamp 1717166647
transform -1 0 3249 0 1 397
box -1519 -797 1519 797
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM8
timestamp 1717166647
transform -1 0 1986 0 1 -3670
box -278 -758 278 758
<< labels >>
flabel metal3 4883 4344 5083 4544 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 -280 2855 -80 3055 0 FreeSans 256 0 0 0 vinn
port 3 nsew
flabel metal2 5026 -3705 5226 -3505 0 FreeSans 256 0 0 0 oneg
port 5 nsew
flabel metal2 5026 -3433 5226 -3233 0 FreeSans 256 0 0 0 opos
port 6 nsew
flabel metal3 -230 -4403 -30 -4203 0 FreeSans 256 0 0 0 avss
port 7 nsew
flabel metal1 -274 1237 -74 1437 0 FreeSans 256 0 0 0 vinp
port 4 nsew
flabel metal1 7630 -158 7830 42 0 FreeSans 256 0 0 0 clka
port 2 nsew
flabel metal1 7642 1464 7842 1664 0 FreeSans 256 0 0 0 enab
port 1 nsew
flabel metal2 6471 -577 6906 -488 0 FreeSans 800 0 0 0 dvdd
port 8 nsew
flabel metal2 7105 -562 7540 -473 0 FreeSans 800 0 0 0 dvss
port 9 nsew
<< end >>
