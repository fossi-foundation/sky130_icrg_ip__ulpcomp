magic
tech sky130A
magscale 1 2
timestamp 1717166647
<< nwell >>
rect -487 -5415 487 5415
<< mvpmos >>
rect -229 118 -29 5118
rect 29 118 229 5118
rect -229 -5118 -29 -118
rect 29 -5118 229 -118
<< mvpdiff >>
rect -287 5106 -229 5118
rect -287 130 -275 5106
rect -241 130 -229 5106
rect -287 118 -229 130
rect -29 5106 29 5118
rect -29 130 -17 5106
rect 17 130 29 5106
rect -29 118 29 130
rect 229 5106 287 5118
rect 229 130 241 5106
rect 275 130 287 5106
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -5106 -275 -130
rect -241 -5106 -229 -130
rect -287 -5118 -229 -5106
rect -29 -130 29 -118
rect -29 -5106 -17 -130
rect 17 -5106 29 -130
rect -29 -5118 29 -5106
rect 229 -130 287 -118
rect 229 -5106 241 -130
rect 275 -5106 287 -130
rect 229 -5118 287 -5106
<< mvpdiffc >>
rect -275 130 -241 5106
rect -17 130 17 5106
rect 241 130 275 5106
rect -275 -5106 -241 -130
rect -17 -5106 17 -130
rect 241 -5106 275 -130
<< mvnsubdiff >>
rect -421 5337 421 5349
rect -421 5303 -313 5337
rect 313 5303 421 5337
rect -421 5291 421 5303
rect -421 5241 -363 5291
rect -421 -5241 -409 5241
rect -375 -5241 -363 5241
rect 363 5241 421 5291
rect -421 -5291 -363 -5241
rect 363 -5241 375 5241
rect 409 -5241 421 5241
rect 363 -5291 421 -5241
rect -421 -5303 421 -5291
rect -421 -5337 -313 -5303
rect 313 -5337 421 -5303
rect -421 -5349 421 -5337
<< mvnsubdiffcont >>
rect -313 5303 313 5337
rect -409 -5241 -375 5241
rect 375 -5241 409 5241
rect -313 -5337 313 -5303
<< poly >>
rect -229 5199 -29 5215
rect -229 5165 -213 5199
rect -45 5165 -29 5199
rect -229 5118 -29 5165
rect 29 5199 229 5215
rect 29 5165 45 5199
rect 213 5165 229 5199
rect 29 5118 229 5165
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -5165 -29 -5118
rect -229 -5199 -213 -5165
rect -45 -5199 -29 -5165
rect -229 -5215 -29 -5199
rect 29 -5165 229 -5118
rect 29 -5199 45 -5165
rect 213 -5199 229 -5165
rect 29 -5215 229 -5199
<< polycont >>
rect -213 5165 -45 5199
rect 45 5165 213 5199
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -5199 -45 -5165
rect 45 -5199 213 -5165
<< locali >>
rect -409 5303 -313 5337
rect 313 5303 409 5337
rect -409 5241 -375 5303
rect 375 5241 409 5303
rect -229 5165 -213 5199
rect -45 5165 -29 5199
rect 29 5165 45 5199
rect 213 5165 229 5199
rect -275 5106 -241 5122
rect -275 114 -241 130
rect -17 5106 17 5122
rect -17 114 17 130
rect 241 5106 275 5122
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -5122 -241 -5106
rect -17 -130 17 -114
rect -17 -5122 17 -5106
rect 241 -130 275 -114
rect 241 -5122 275 -5106
rect -229 -5199 -213 -5165
rect -45 -5199 -29 -5165
rect 29 -5199 45 -5165
rect 213 -5199 229 -5165
rect -409 -5303 -375 -5241
rect 375 -5303 409 -5241
rect -409 -5337 -313 -5303
rect 313 -5337 409 -5303
<< viali >>
rect -213 5165 -45 5199
rect 45 5165 213 5199
rect -275 130 -241 5106
rect -17 130 17 5106
rect 241 130 275 5106
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -5106 -241 -130
rect -17 -5106 17 -130
rect 241 -5106 275 -130
rect -213 -5199 -45 -5165
rect 45 -5199 213 -5165
<< metal1 >>
rect -225 5199 -33 5205
rect -225 5165 -213 5199
rect -45 5165 -33 5199
rect -225 5159 -33 5165
rect 33 5199 225 5205
rect 33 5165 45 5199
rect 213 5165 225 5199
rect 33 5159 225 5165
rect -281 5106 -235 5118
rect -281 130 -275 5106
rect -241 130 -235 5106
rect -281 118 -235 130
rect -23 5106 23 5118
rect -23 130 -17 5106
rect 17 130 23 5106
rect -23 118 23 130
rect 235 5106 281 5118
rect 235 130 241 5106
rect 275 130 281 5106
rect 235 118 281 130
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -130 -235 -118
rect -281 -5106 -275 -130
rect -241 -5106 -235 -130
rect -281 -5118 -235 -5106
rect -23 -130 23 -118
rect -23 -5106 -17 -130
rect 17 -5106 23 -130
rect -23 -5118 23 -5106
rect 235 -130 281 -118
rect 235 -5106 241 -130
rect 275 -5106 281 -130
rect 235 -5118 281 -5106
rect -225 -5165 -33 -5159
rect -225 -5199 -213 -5165
rect -45 -5199 -33 -5165
rect -225 -5205 -33 -5199
rect 33 -5165 225 -5159
rect 33 -5199 45 -5165
rect 213 -5199 225 -5165
rect 33 -5205 225 -5199
<< properties >>
string FIXED_BBOX -392 -5320 392 5320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 25.0 l 1.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
