** sch_path: /home/ttuser/chipalooza2024/sky130_icrg_ip__ulpcomp/cace/tb_static_current.sch
**.subckt tb_static_current
V3 ena GND {ena}*{dvdd}
avdd avdd GND {avdd}
dvdd dvdd GND {dvdd}
avss avss GND {avss}
dvss dvss GND {dvss}
Vcm vinn GND VOL=' {Vcm} '
XC1 vout GND sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=3 m=3
x1 dvdd avdd ena vinp vinn vout net1 avss dvss sky130_icrg_ip__ulpcomp
Vdiff vinp vinn {Vdiff}
**** begin user architecture code


.lib /home/ttuser/pdk/sky130A/libs.tech/combined/sky130.lib.spice {corner}
.option TEMP={temperature}


.control
op
set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -I(dvdd)
quit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
