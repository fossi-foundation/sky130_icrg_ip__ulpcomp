* NGSPICE file created from sky130_icrg_ip__ulpcomp2.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_PVEW3M a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_XPB8Y6 a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt Stage0_clk_inv dvddb clka clk clkb dvss
XXM6 dvss clkb dvss clk sky130_fd_pr__nfet_01v8_PVEW3M
XXM8 clkb clka dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
XXM21 dvss clka dvss clkb sky130_fd_pr__nfet_01v8_PVEW3M
XXM22 clk clkb dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.12188 ps=1.075 w=0.75 l=0.5
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X12 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.12188 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGL9FS a_29_n597# a_n287_n500# a_n229_n597# a_287_n597#
+ a_229_n500# w_n745_n797# a_n545_n500# a_n487_n597# a_n29_n500# a_487_n500#
X0 a_487_n500# a_287_n597# a_229_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_229_n500# a_29_n597# a_n29_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n597# a_n287_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E2TVSU a_1261_n500# a_n1319_n500# a_29_n597#
+ a_n287_n500# a_n1061_n500# a_n745_n597# a_803_n597# a_745_n500# a_n229_n597# a_287_n597#
+ a_n1003_n597# a_229_n500# w_n1519_n797# a_n545_n500# a_1061_n597# a_1003_n500# a_n487_n597#
+ a_n1261_n597# a_n29_n500# a_545_n597# a_487_n500# a_n803_n500#
X0 a_n1061_n500# a_n1261_n597# a_n1319_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X1 a_1003_n500# a_803_n597# a_745_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_487_n500# a_287_n597# a_229_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_745_n500# a_545_n597# a_487_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1261_n500# a_1061_n597# a_1003_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_229_n500# a_29_n597# a_n29_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n29_n500# a_n229_n597# a_n287_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n500# a_n745_n597# a_n803_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_n287_n500# a_n487_n597# a_n545_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n803_n500# a_n1003_n597# a_n1061_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_03v3_nvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt Stage1 enab clka vinn vinp oneg opos avss avdd w_608_n4673# dvdd dvss
Xx1 clka dvdd dvss dvss avdd avdd x1/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xx2 enab dvdd dvss dvss avdd avdd x2/X sky130_fd_sc_hvl__lsbuflv2hv_1
XXM3_2 vinp oneg vinp vinp oneg li_n3_908# li_n3_908# vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM1_1 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM1_2 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM5 opos w_608_n4673# w_608_n4673# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM6_1 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM6_2 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM8 oneg w_608_n4673# w_608_n4673# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM4_2 avss avss w_608_n4673# w_608_n4673# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_0 vinp oneg vinp vinp oneg li_n3_908# li_n3_908#
+ vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_1 vinn opos vinn vinn opos li_n3_908# li_n3_908#
+ vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM2_2 vinn opos vinn vinn opos li_n3_908# li_n3_908# vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__nfet_03v3_nvt_FJGQ2Y_0 avss avss w_608_n4673# w_608_n4673# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8_hvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_03v3_nvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_3HY9VM w_n296_n419# a_n100_n297# a_100_n200# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n296_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt Stage2_latch dvdd enab dvddb clkb vout oneg opos dvss
XXM12 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM15 dvss dvss m2_1568_n2406# clkb sky130_fd_pr__nfet_03v3_nvt_WSEQJ8
XXM18 dvss dvss vout m1_683_n2348# sky130_fd_pr__nfet_01v8_PVEW3M
XXM19 dvddb m1_683_n2348# dvddb vout sky130_fd_pr__pfet_01v8_3HY9VM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_0 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM1 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_1 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_3 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_2 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM2 dvss m1_1866_n2368# m1_683_n2348# opos sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_4 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM3 dvss m2_1568_n2406# m1_1866_n2368# m2_1331_n391# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_5 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM4 dvss m1_2747_n2368# m2_1331_n391# oneg sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM5 dvss m2_1568_n2406# m1_2747_n2368# m1_683_n2348# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM10 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM11 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
.ends

.subckt Stage0_ena_inv dvdd ena enab dvss
XXM25 ena enab dvdd dvdd sky130_fd_pr__pfet_01v8_XPB8Y6
XXM24 dvss enab dvss ena sky130_fd_pr__nfet_01v8_PVEW3M
.ends

.subckt sky130_icrg_ip__ulpcomp2 avdd ena vout vinn vinp dvss avss clk dvdd
Xx1 x3/dvddb x2/clka clk x3/clkb dvss Stage0_clk_inv
Xx2 x4/enab x2/clka vinn vinp x3/oneg x3/opos avss avdd w_288_n7721# dvdd dvss Stage1
Xx3 dvdd x4/enab x3/dvddb x3/clkb vout x3/oneg x3/opos dvss Stage2_latch
Xx4 dvdd ena x4/enab dvss Stage0_ena_inv
.ends

