magic
tech sky130A
magscale 1 2
timestamp 1747754763
<< psubdiff >>
rect -576 1530 -516 1564
rect 8444 1530 8504 1564
rect -576 1504 -542 1530
rect 8470 1504 8504 1530
rect -344 -5279 -320 -5165
rect 4455 -5279 4479 -5165
rect -576 -8122 -542 -8096
rect 8470 -8122 8504 -8096
rect -576 -8156 -516 -8122
rect 8444 -8156 8504 -8122
<< psubdiffcont >>
rect -516 1530 8444 1564
rect -576 -8096 -542 1504
rect -320 -5279 4455 -5165
rect 8470 -8096 8504 1504
rect -516 -8156 8444 -8122
<< locali >>
rect -576 1553 -516 1564
rect 8444 1553 8504 1564
rect -576 1511 -549 1553
rect 8469 1511 8504 1553
rect -576 1504 8504 1511
rect -542 1433 8470 1504
rect -542 -5051 -490 1433
rect -542 -5165 4607 -5051
rect -542 -5279 -320 -5165
rect 4455 -5279 4607 -5165
rect -542 -5378 4607 -5279
rect -542 -8069 -490 -5378
rect 8430 -8069 8470 1433
rect -542 -8086 8470 -8069
rect 8466 -8096 8470 -8086
rect -576 -8133 -548 -8096
rect 8466 -8133 8504 -8096
rect -576 -8156 -516 -8133
rect 8444 -8156 8504 -8133
<< viali >>
rect -549 1530 -516 1553
rect -516 1530 8444 1553
rect 8444 1530 8469 1553
rect -549 1511 8469 1530
rect -548 -8096 -542 -8086
rect -542 -8096 8466 -8086
rect -548 -8122 8466 -8096
rect -548 -8133 -516 -8122
rect -516 -8133 8444 -8122
rect 8444 -8133 8466 -8122
<< metal1 >>
rect -576 1553 8504 1565
rect -576 1511 -549 1553
rect 8469 1511 8504 1553
rect -576 1490 8504 1511
rect 6262 1411 6451 1490
rect 7354 1462 8225 1490
rect 7698 1415 7887 1462
rect 6580 818 6757 862
rect 6011 735 6122 773
rect -600 -193 -400 7
rect 6011 -76 6049 735
rect 6713 4 6757 818
rect 8113 726 8265 926
rect 6713 -40 8242 4
rect 6011 -114 7750 -76
rect 7713 -1492 7750 -114
rect 8090 -216 8242 -40
rect 7466 -1530 7960 -1492
rect -594 -1811 -394 -1611
rect 7678 -3128 7716 -3052
rect 7466 -3166 7716 -3128
rect 7463 -3679 7713 -3644
rect 7463 -3897 7498 -3679
rect 7925 -3744 7960 -1530
rect 7750 -3779 7960 -3744
rect 7750 -3891 7785 -3779
rect 7754 -3892 7785 -3891
rect 8264 -6897 8464 -6697
rect 5373 -8070 5573 -7298
rect 7320 -8070 7520 -7306
rect -568 -8086 8495 -8070
rect -568 -8133 -548 -8086
rect 8466 -8133 8495 -8086
rect -568 -8148 8495 -8133
<< metal2 >>
rect 6402 1268 8239 1474
rect 6150 -194 6585 231
rect 6325 -195 6585 -194
rect 6783 -250 6990 1268
rect 7141 730 7490 769
rect 7141 -81 7180 730
rect 7821 682 7860 763
rect 7229 643 7860 682
rect 7229 -9 7268 643
rect 7229 -48 7813 -9
rect 7141 -120 7718 -81
rect 6151 -2057 6586 -2026
rect 7679 -3039 7718 -120
rect 7774 -3211 7813 -48
rect 7679 -3250 7813 -3211
rect 7679 -3484 7718 -3250
rect 7880 -3318 8039 57
rect 7826 -3477 8039 -3318
rect 6784 -3540 7221 -3529
rect 6784 -3662 6799 -3540
rect 7205 -3662 7221 -3540
rect 6784 -3679 7221 -3662
rect 7826 -4405 7985 -3477
rect 8104 -3596 8334 -3578
rect 8104 -3871 8121 -3596
rect 8309 -3871 8334 -3596
rect 8104 -3907 8334 -3871
rect 7304 -7195 7533 -7187
rect 7304 -7379 7313 -7195
rect 7523 -7379 7533 -7195
rect 7304 -7386 7533 -7379
rect 7846 -7387 8222 -7187
<< via2 >>
rect 6162 -3340 6571 -3212
rect 6799 -3662 7205 -3540
rect 8121 -3871 8309 -3596
rect 7313 -7379 7523 -7195
<< metal3 >>
rect 4475 1495 4904 1566
rect 4475 1071 4903 1495
rect 6150 -3212 8329 -3201
rect 6150 -3340 6162 -3212
rect 6571 -3340 8329 -3212
rect 6150 -3388 8329 -3340
rect 6784 -3540 7581 -3526
rect 6784 -3662 6799 -3540
rect 7205 -3662 7581 -3540
rect 6784 -3710 7581 -3662
rect -624 -7460 -196 -6947
rect 7304 -7187 7581 -3710
rect 8105 -3596 8329 -3388
rect 8105 -3871 8121 -3596
rect 8309 -3871 8329 -3596
rect 8105 -3886 8329 -3871
rect 7304 -7195 8222 -7187
rect 7304 -7379 7313 -7195
rect 7523 -7379 8222 -7195
rect 7304 -7387 8222 -7379
rect -625 -8146 -196 -7460
use pa_via_short  pa_via_short_0
timestamp 1717168741
transform -1 0 12673 0 1 -1794
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_1
timestamp 1717168741
transform -1 0 12673 0 1 -1279
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_2
timestamp 1717168741
transform -1 0 12831 0 1 2609
box 4944 -1889 5010 -1683
use pa_via_short  pa_via_short_22
timestamp 1717168741
transform -1 0 12455 0 1 2605
box 4944 -1889 5010 -1683
use Stage0_clk_inv  x1
timestamp 1717191815
transform -1 0 8551 0 -1 215
box 321 -1284 1222 196
use Stage1  x2
timestamp 1747754759
transform 1 0 -320 0 1 -3048
box -305 -4988 7963 4550
use Stage2_latch  x3
timestamp 1747754763
transform -1 0 8763 0 1 -4587
box 300 -2867 4057 739
use Stage0_ena_inv  x4
timestamp 1717183580
transform -1 0 6992 0 -1 169
box 379 -1306 885 152
<< labels >>
flabel metal3 8022 -7387 8222 -7187 0 FreeSans 960 0 0 0 dvss
port 7 nsew
flabel metal1 8113 726 8265 926 0 FreeSans 256 0 0 0 clk
port 9 nsew
flabel metal3 4563 1296 4763 1494 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 8090 -216 8242 -16 0 FreeSans 256 180 0 0 ena
port 2 nsew
flabel metal3 8105 -3596 8329 -3201 0 FreeSans 1120 90 0 0 dvdd
port 10 nsew
flabel metal1 8264 -6897 8464 -6697 0 FreeSans 256 0 0 0 vout
port 3 nsew
flabel metal1 -600 -193 -400 7 0 FreeSans 256 0 0 0 vinn
port 4 nsew
flabel metal1 -594 -1811 -394 -1611 0 FreeSans 256 0 0 0 vinp
port 5 nsew
flabel metal3 -549 -7450 -349 -7250 0 FreeSans 256 0 0 0 avss
port 8 nsew
<< end >>
