** sch_path: /home/ttuser/chipalooza2024/sky130_icrg_ip__ulpcomp/cace/tb_dynamic_current.sch
**.subckt tb_dynamic_current
V3 ena GND Pulse(0 {ena}*1.8 0 0.1n 0.1n 0.5n 1n)
avdd avdd GND {avdd}
dvdd dvdd GND {dvdd}
avss avss GND {avss}
dvss dvss GND {dvss}
E1 vinn GND VOL=' DC 0 sin(0 {Vdiff} {frequency2} 0 0) '
E2 vinp GND VOL=' DC 0 sin(0 {Vdiff} {frequency1} 0 0) '
XC1 vout GND sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=3 m=3
x1 dvdd avdd ena vinp vinn vout net1 avss dvss sky130_icrg_ip__ulpcomp
**** begin user architecture code


.lib /home/ttuser/pdk/sky130A/libs.tech/combined/sky130.lib.spice {corner}
.option TEMP={temperature}


.control
tran [1.0 / {frequency1} / 100] [1 / {frequency1}]
set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -I(dvdd)
quit
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
